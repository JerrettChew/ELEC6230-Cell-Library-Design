magic
tech tsmc180
timestamp 1733141978
<< nwell >>
rect 0 637 186 1176
<< polysilicon >>
rect 66 1110 75 1121
rect 102 1110 111 1121
rect 141 1110 150 1121
rect 66 1005 75 1021
rect 102 1005 111 1021
rect 141 977 150 1021
rect 66 902 75 916
rect 102 902 111 916
rect 66 206 75 877
rect 102 206 111 877
rect 141 239 150 956
rect 66 121 75 157
rect 102 121 111 157
rect 141 121 150 218
rect 66 61 75 72
rect 102 61 111 72
rect 141 61 150 72
<< ndiffusion >>
rect 63 157 66 206
rect 75 157 78 206
rect 99 157 102 206
rect 111 157 114 206
rect 63 72 66 121
rect 75 72 102 121
rect 111 72 114 121
rect 135 72 141 121
rect 150 72 153 121
<< pdiffusion >>
rect 63 1021 66 1110
rect 75 1021 78 1110
rect 99 1021 102 1110
rect 111 1021 114 1110
rect 135 1021 141 1110
rect 150 1021 154 1110
rect 63 916 66 1005
rect 75 916 102 1005
rect 111 916 115 1005
<< pohmic >>
rect 0 15 2 36
rect 23 15 33 36
rect 54 15 66 36
rect 87 15 99 36
rect 120 15 132 36
rect 153 15 162 36
rect 183 15 186 36
<< nohmic >>
rect 0 1146 2 1167
rect 23 1146 33 1167
rect 54 1146 66 1167
rect 87 1146 99 1167
rect 120 1146 132 1167
rect 153 1146 162 1167
rect 183 1146 186 1167
<< ntransistor >>
rect 66 157 75 206
rect 102 157 111 206
rect 66 72 75 121
rect 102 72 111 121
rect 141 72 150 121
<< ptransistor >>
rect 66 1021 75 1110
rect 102 1021 111 1110
rect 141 1021 150 1110
rect 66 916 75 1005
rect 102 916 111 1005
<< polycontact >>
rect 141 956 162 977
rect 54 877 80 902
rect 99 877 123 902
rect 129 218 150 239
<< ndiffcontact >>
rect 42 157 63 206
rect 78 157 99 206
rect 114 157 135 206
rect 42 72 63 121
rect 114 72 135 121
rect 153 72 174 121
<< pdiffcontact >>
rect 42 1021 63 1110
rect 78 1021 99 1110
rect 114 1021 135 1110
rect 154 1021 175 1110
rect 42 916 63 1005
rect 115 916 136 1005
<< psubstratetap >>
rect 2 15 23 36
rect 33 15 54 36
rect 66 15 87 36
rect 99 15 120 36
rect 132 15 153 36
rect 162 15 183 36
<< nsubstratetap >>
rect 2 1146 23 1167
rect 33 1146 54 1167
rect 66 1146 87 1167
rect 99 1146 120 1167
rect 132 1146 153 1167
rect 162 1146 183 1167
<< metal1 >>
rect 0 1167 186 1176
rect 0 1146 2 1167
rect 23 1146 33 1167
rect 54 1146 66 1167
rect 87 1146 99 1167
rect 120 1146 132 1167
rect 153 1146 162 1167
rect 183 1146 186 1167
rect 6 1005 30 1146
rect 42 1122 135 1134
rect 42 1110 63 1122
rect 114 1110 135 1122
rect 78 1005 99 1021
rect 6 916 42 1005
rect 63 916 99 1005
rect 136 956 141 977
rect 0 546 186 558
rect 0 517 186 529
rect 0 488 186 500
rect 0 459 186 471
rect 0 430 186 442
rect 78 218 129 230
rect 78 206 99 218
rect 42 145 63 157
rect 114 145 135 157
rect 6 133 135 145
rect 6 36 30 133
rect 114 121 135 133
rect 42 60 63 72
rect 153 60 174 72
rect 42 48 174 60
rect 0 15 2 36
rect 23 15 33 36
rect 54 15 66 36
rect 87 15 99 36
rect 120 15 132 36
rect 153 15 162 36
rect 183 15 186 36
rect 0 6 186 15
<< m2contact >>
rect 160 1081 175 1100
rect 175 1081 179 1100
rect 54 877 80 902
rect 99 877 123 902
rect 160 100 174 119
rect 174 100 179 119
<< metal2 >>
rect 66 902 80 1182
rect 66 0 80 877
rect 99 902 113 1182
rect 165 1100 179 1182
rect 99 0 113 877
rect 165 119 179 1081
rect 165 0 179 100
<< labels >>
rlabel polysilicon 106 61 106 61 1 B
rlabel polysilicon 70 61 70 61 1 A
rlabel polysilicon 145 61 145 61 1 n1
rlabel metal2 165 0 179 0 1 Y
rlabel metal2 99 0 113 0 1 B
rlabel metal2 66 0 80 0 1 A
rlabel metal1 0 6 0 36 3 GND!
rlabel metal1 186 6 186 36 7 GND!
rlabel metal2 99 1182 113 1182 5 B
rlabel metal2 165 1182 179 1182 5 Y
rlabel metal2 66 1182 80 1182 5 A
rlabel polysilicon 145 1121 145 1121 1 n1
rlabel polysilicon 71 1121 71 1121 1 A
rlabel polysilicon 106 1121 106 1121 1 B
rlabel metal1 186 1146 186 1176 7 Vdd!
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 430 0 442 3 nReset
rlabel metal1 186 488 186 500 7 Test
rlabel metal1 186 459 186 471 7 Clock
rlabel metal1 186 430 186 442 7 nReset
rlabel metal1 0 546 0 558 3 Scan
rlabel metal1 186 546 186 558 7 Scan
rlabel metal1 186 517 186 529 7 ScanReturn
rlabel metal1 0 517 0 529 3 ScanReturn
<< end >>
