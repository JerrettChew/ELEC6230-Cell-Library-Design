magic
tech tsmc180
timestamp 1732895094
<< nwell >>
rect 0 637 301 1176
<< polysilicon >>
rect 73 1119 82 1130
rect 109 1119 118 1130
rect 147 1119 156 1130
rect 73 994 82 1030
rect 109 994 118 1030
rect 147 994 156 1030
rect 185 994 194 1130
rect 261 1051 270 1130
rect 73 851 82 905
rect 109 851 118 905
rect 73 726 82 762
rect 109 726 118 762
rect 147 726 156 905
rect 185 851 194 905
rect 261 851 270 1030
rect 73 625 82 637
rect 73 385 82 604
rect 109 591 118 637
rect 147 591 156 637
rect 185 625 194 762
rect 190 604 194 625
rect 109 385 118 570
rect 147 385 156 570
rect 185 418 194 604
rect 190 397 194 418
rect 73 300 82 336
rect 109 300 118 336
rect 73 197 82 251
rect 109 197 118 251
rect 147 197 156 336
rect 185 300 194 397
rect 261 300 270 762
rect 185 197 194 251
rect 73 112 82 148
rect 109 112 118 148
rect 147 112 156 148
rect 73 52 82 63
rect 109 52 118 63
rect 147 52 156 63
rect 185 52 194 148
rect 261 112 270 251
rect 261 52 270 91
<< ndiffusion >>
rect 70 336 73 385
rect 82 336 109 385
rect 118 336 121 385
rect 142 336 147 385
rect 156 336 159 385
rect 70 251 73 300
rect 82 251 85 300
rect 106 251 109 300
rect 118 251 121 300
rect 182 251 185 300
rect 194 251 202 300
rect 258 251 261 300
rect 270 251 273 300
rect 70 148 73 197
rect 82 148 85 197
rect 106 148 109 197
rect 118 148 121 197
rect 142 148 147 197
rect 156 148 159 197
rect 180 148 185 197
rect 194 148 202 197
rect 70 63 73 112
rect 82 63 109 112
rect 118 63 147 112
rect 156 63 159 112
<< pdiffusion >>
rect 70 1030 73 1119
rect 82 1030 109 1119
rect 118 1030 147 1119
rect 156 1030 159 1119
rect 70 905 73 994
rect 82 905 85 994
rect 106 905 109 994
rect 118 905 121 994
rect 142 905 147 994
rect 156 905 159 994
rect 180 905 185 994
rect 194 905 202 994
rect 70 762 73 851
rect 82 762 85 851
rect 106 762 109 851
rect 118 762 121 851
rect 182 762 185 851
rect 194 762 202 851
rect 258 762 261 851
rect 270 762 273 851
rect 70 637 73 726
rect 82 637 109 726
rect 118 637 121 726
rect 142 637 147 726
rect 156 637 159 726
<< pohmic >>
rect 0 15 33 36
rect 54 15 66 36
rect 87 15 99 36
rect 120 15 132 36
rect 153 15 165 36
rect 186 15 198 36
rect 219 15 231 36
rect 252 15 264 36
rect 285 15 301 36
<< nohmic >>
rect 0 1146 33 1167
rect 54 1146 66 1167
rect 87 1146 99 1167
rect 120 1146 132 1167
rect 153 1146 165 1167
rect 186 1146 198 1167
rect 219 1146 231 1167
rect 252 1146 264 1167
rect 285 1146 301 1167
<< ntransistor >>
rect 73 336 82 385
rect 109 336 118 385
rect 147 336 156 385
rect 73 251 82 300
rect 109 251 118 300
rect 185 251 194 300
rect 261 251 270 300
rect 73 148 82 197
rect 109 148 118 197
rect 147 148 156 197
rect 185 148 194 197
rect 73 63 82 112
rect 109 63 118 112
rect 147 63 156 112
<< ptransistor >>
rect 73 1030 82 1119
rect 109 1030 118 1119
rect 147 1030 156 1119
rect 73 905 82 994
rect 109 905 118 994
rect 147 905 156 994
rect 185 905 194 994
rect 73 762 82 851
rect 109 762 118 851
rect 185 762 194 851
rect 261 762 270 851
rect 73 637 82 726
rect 109 637 118 726
rect 147 637 156 726
<< polycontact >>
rect 249 1030 270 1051
rect 67 604 88 625
rect 169 604 190 625
rect 103 570 124 591
rect 141 570 162 591
rect 169 397 190 418
rect 249 91 270 112
<< ndiffcontact >>
rect 49 336 70 385
rect 121 336 142 385
rect 159 336 180 385
rect 49 251 70 300
rect 85 251 106 300
rect 121 251 142 300
rect 161 251 182 300
rect 202 251 223 300
rect 237 251 258 300
rect 273 251 294 300
rect 49 148 70 197
rect 85 148 106 197
rect 121 148 142 197
rect 159 148 180 197
rect 202 148 223 197
rect 49 63 70 112
rect 159 63 180 112
<< pdiffcontact >>
rect 49 1030 70 1119
rect 159 1030 180 1119
rect 49 905 70 994
rect 85 905 106 994
rect 121 905 142 994
rect 159 905 180 994
rect 202 905 223 994
rect 49 762 70 851
rect 85 762 106 851
rect 121 762 142 851
rect 161 762 182 851
rect 202 762 223 851
rect 237 762 258 851
rect 273 762 294 851
rect 49 637 70 726
rect 121 637 142 726
rect 159 637 180 726
<< psubstratetap >>
rect 33 15 54 36
rect 66 15 87 36
rect 99 15 120 36
rect 132 15 153 36
rect 165 15 186 36
rect 198 15 219 36
rect 231 15 252 36
rect 264 15 285 36
<< nsubstratetap >>
rect 33 1146 54 1167
rect 66 1146 87 1167
rect 99 1146 120 1167
rect 132 1146 153 1167
rect 165 1146 186 1167
rect 198 1146 219 1167
rect 231 1146 252 1167
rect 264 1146 285 1167
<< metal1 >>
rect 0 1167 301 1176
rect 0 1146 33 1167
rect 54 1146 66 1167
rect 87 1146 99 1167
rect 120 1146 132 1167
rect 153 1146 165 1167
rect 186 1146 198 1167
rect 219 1146 231 1167
rect 252 1146 264 1167
rect 285 1146 301 1167
rect 7 893 37 1146
rect 180 1030 249 1042
rect 49 1018 70 1030
rect 49 1006 180 1018
rect 85 994 106 1006
rect 159 994 180 1006
rect 211 994 223 1030
rect 49 893 70 905
rect 121 893 142 905
rect 7 863 294 893
rect 85 851 106 863
rect 161 851 182 863
rect 237 851 258 863
rect 49 750 70 762
rect 121 750 142 762
rect 49 738 180 750
rect 49 726 70 738
rect 159 726 180 738
rect 125 621 137 637
rect 125 609 169 621
rect 211 623 223 762
rect 282 623 294 762
rect 211 611 229 623
rect 281 611 294 623
rect 162 572 163 591
rect 0 546 301 558
rect 0 517 301 529
rect 0 488 301 500
rect 0 459 301 471
rect 0 430 301 442
rect 125 402 169 414
rect 125 385 137 402
rect 211 399 229 411
rect 281 399 294 411
rect 49 324 70 336
rect 161 324 180 336
rect 49 312 180 324
rect 49 300 70 312
rect 121 300 142 312
rect 211 300 223 399
rect 282 300 294 399
rect 85 239 106 251
rect 161 239 180 251
rect 237 239 258 251
rect 7 209 294 239
rect 7 36 37 209
rect 49 197 70 209
rect 121 197 142 209
rect 85 136 106 148
rect 159 136 180 148
rect 49 124 180 136
rect 49 112 70 124
rect 211 112 223 148
rect 180 100 249 112
rect 0 15 33 36
rect 54 15 66 36
rect 87 15 99 36
rect 120 15 132 36
rect 153 15 165 36
rect 186 15 198 36
rect 219 15 231 36
rect 252 15 264 36
rect 285 15 301 36
rect 0 6 301 15
<< m2contact >>
rect 61 606 67 625
rect 67 606 80 625
rect 229 604 248 623
rect 262 604 281 623
rect 97 572 103 591
rect 103 572 116 591
rect 163 572 182 591
rect 229 399 248 418
rect 262 399 281 418
<< metal2 >>
rect 66 625 80 1182
rect 66 0 80 606
rect 99 591 113 1182
rect 165 591 179 1182
rect 231 623 245 1182
rect 264 623 278 1182
rect 99 0 113 572
rect 165 0 179 572
rect 231 418 245 604
rect 264 418 278 604
rect 231 0 245 399
rect 264 0 278 399
<< labels >>
rlabel polysilicon 190 1130 190 1130 1 D
rlabel polysilicon 190 52 190 52 1 D
rlabel polysilicon 263 1130 263 1130 1 Y
rlabel polysilicon 263 52 263 52 1 Y
rlabel metal2 264 1182 278 1182 5 S
rlabel metal2 231 1182 245 1182 5 Cout
rlabel metal2 165 1182 179 1182 5 Cin
rlabel metal2 99 1182 113 1182 5 B
rlabel metal2 66 1182 80 1182 5 A
rlabel metal2 66 0 80 0 1 A
rlabel metal2 99 0 113 0 1 B
rlabel metal2 165 0 179 0 1 Cin
rlabel metal2 231 0 245 0 1 Cout
rlabel metal2 264 0 278 0 1 S
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel metal1 301 1146 301 1176 7 Vdd!
rlabel metal1 0 6 0 36 3 GND!
rlabel metal1 301 6 301 36 7 GND!
rlabel metal1 0 546 0 558 3 Scan
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 430 0 442 3 nReset
rlabel metal1 301 546 301 558 7 Scan
rlabel metal1 301 517 301 529 7 ScanReturn
rlabel metal1 301 488 301 500 7 Test
rlabel metal1 301 459 301 471 7 Clock
rlabel metal1 301 430 301 442 7 nReset
<< end >>
