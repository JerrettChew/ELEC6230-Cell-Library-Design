magic
tech tsmc180
timestamp 1733141177
<< nwell >>
rect 0 637 398 1176
<< polysilicon >>
rect 54 915 63 1141
rect 92 1053 101 1141
rect 130 1110 139 1141
rect 130 1089 134 1110
rect 130 1053 139 1089
rect 168 1053 177 1141
rect 204 1053 213 1141
rect 54 757 63 826
rect 92 757 101 964
rect 130 915 139 964
rect 168 915 177 964
rect 204 915 213 964
rect 54 352 63 668
rect 92 475 101 668
rect 92 352 101 454
rect 54 245 63 303
rect 54 41 63 196
rect 92 147 101 303
rect 130 245 139 826
rect 168 790 177 826
rect 173 769 177 790
rect 168 757 177 769
rect 204 757 213 826
rect 242 814 251 1141
rect 280 1053 289 1141
rect 320 1134 329 1141
rect 320 1053 329 1113
rect 242 757 251 793
rect 168 352 177 668
rect 204 446 213 668
rect 242 562 251 668
rect 280 593 289 964
rect 320 915 329 964
rect 358 915 367 1141
rect 204 352 213 425
rect 242 352 251 541
rect 168 278 177 303
rect 168 245 177 257
rect 204 245 213 303
rect 242 278 251 303
rect 130 147 139 196
rect 168 147 177 196
rect 204 147 213 196
rect 92 41 101 98
rect 130 93 139 98
rect 130 41 139 72
rect 168 41 177 98
rect 204 41 213 98
rect 242 41 251 257
rect 280 147 289 572
rect 320 245 329 826
rect 358 757 367 826
rect 358 591 367 668
rect 358 352 367 570
rect 358 245 367 303
rect 320 147 329 196
rect 280 41 289 98
rect 320 69 329 98
rect 320 41 329 48
rect 358 41 367 196
<< ndiffusion >>
rect 51 303 54 352
rect 63 303 92 352
rect 101 303 104 352
rect 165 303 168 352
rect 177 303 204 352
rect 213 303 242 352
rect 251 303 254 352
rect 127 196 130 245
rect 139 196 168 245
rect 177 196 204 245
rect 213 196 216 245
rect 89 98 92 147
rect 101 98 130 147
rect 139 98 168 147
rect 177 98 204 147
rect 213 98 216 147
rect 317 196 320 245
rect 329 196 358 245
rect 367 196 370 245
rect 277 98 280 147
rect 289 98 320 147
rect 329 98 332 147
<< pdiffusion >>
rect 89 964 92 1053
rect 101 964 104 1053
rect 125 964 130 1053
rect 139 964 142 1053
rect 163 964 168 1053
rect 177 964 180 1053
rect 201 964 204 1053
rect 213 964 216 1053
rect 127 826 130 915
rect 139 826 142 915
rect 163 826 168 915
rect 177 826 180 915
rect 201 826 204 915
rect 213 826 216 915
rect 51 668 54 757
rect 63 668 66 757
rect 87 668 92 757
rect 101 668 104 757
rect 277 964 280 1053
rect 289 964 292 1053
rect 313 964 320 1053
rect 329 964 332 1053
rect 165 668 168 757
rect 177 668 180 757
rect 201 668 204 757
rect 213 668 216 757
rect 237 668 242 757
rect 251 668 254 757
rect 315 826 320 915
rect 329 826 332 915
rect 353 826 358 915
rect 367 826 370 915
<< pohmic >>
rect 0 15 16 36
rect 37 15 68 36
rect 89 15 144 36
rect 165 15 218 36
rect 239 15 292 36
rect 313 15 369 36
rect 390 15 398 36
<< nohmic >>
rect 0 1146 23 1167
rect 44 1146 66 1167
rect 87 1146 144 1167
rect 165 1146 217 1167
rect 238 1146 296 1167
rect 317 1146 368 1167
rect 389 1146 398 1167
<< ntransistor >>
rect 54 303 63 352
rect 92 303 101 352
rect 168 303 177 352
rect 204 303 213 352
rect 242 303 251 352
rect 130 196 139 245
rect 168 196 177 245
rect 204 196 213 245
rect 92 98 101 147
rect 130 98 139 147
rect 168 98 177 147
rect 204 98 213 147
rect 320 196 329 245
rect 358 196 367 245
rect 280 98 289 147
rect 320 98 329 147
<< ptransistor >>
rect 92 964 101 1053
rect 130 964 139 1053
rect 168 964 177 1053
rect 204 964 213 1053
rect 130 826 139 915
rect 168 826 177 915
rect 204 826 213 915
rect 54 668 63 757
rect 92 668 101 757
rect 280 964 289 1053
rect 320 964 329 1053
rect 168 668 177 757
rect 204 668 213 757
rect 242 668 251 757
rect 320 826 329 915
rect 358 826 367 915
<< polycontact >>
rect 134 1089 155 1110
rect 54 826 75 915
rect 92 454 113 475
rect 54 196 75 245
rect 152 769 173 790
rect 308 1113 329 1134
rect 234 793 255 814
rect 268 572 289 593
rect 230 541 251 562
rect 204 425 225 446
rect 156 257 177 278
rect 236 257 257 278
rect 130 72 151 93
rect 346 668 367 757
rect 353 570 374 591
rect 346 303 367 352
rect 308 48 329 69
<< ndiffcontact >>
rect 30 303 51 352
rect 104 303 125 352
rect 144 303 165 352
rect 254 303 275 352
rect 106 196 127 245
rect 216 196 237 245
rect 68 98 89 147
rect 216 98 237 147
rect 294 196 317 245
rect 370 196 391 245
rect 256 98 277 147
rect 332 98 353 147
<< pdiffcontact >>
rect 68 964 89 1053
rect 104 964 125 1053
rect 142 964 163 1053
rect 180 964 201 1053
rect 216 964 237 1053
rect 106 826 127 915
rect 142 826 163 915
rect 180 826 201 915
rect 216 826 237 915
rect 30 668 51 757
rect 66 668 87 757
rect 104 668 125 757
rect 256 964 277 1053
rect 292 964 313 1053
rect 332 964 353 1053
rect 144 668 165 757
rect 180 668 201 757
rect 216 668 237 757
rect 254 668 275 757
rect 294 826 315 915
rect 332 826 353 915
rect 370 826 391 915
<< psubstratetap >>
rect 16 15 37 36
rect 68 15 89 36
rect 144 15 165 36
rect 218 15 239 36
rect 292 15 313 36
rect 369 15 390 36
<< nsubstratetap >>
rect 23 1146 44 1167
rect 66 1146 87 1167
rect 144 1146 165 1167
rect 217 1146 238 1167
rect 296 1146 317 1167
rect 368 1146 389 1167
<< metal1 >>
rect 0 1167 398 1176
rect 0 1146 23 1167
rect 44 1146 66 1167
rect 87 1146 144 1167
rect 165 1146 217 1167
rect 238 1146 296 1167
rect 317 1146 368 1167
rect 389 1146 398 1167
rect 6 952 36 1146
rect 104 1122 308 1134
rect 104 1077 122 1122
rect 155 1089 313 1101
rect 104 1065 201 1077
rect 104 1053 125 1065
rect 180 1053 201 1065
rect 292 1053 313 1089
rect 68 952 89 964
rect 142 952 163 964
rect 216 952 237 964
rect 256 952 277 964
rect 332 952 353 964
rect 6 927 353 952
rect 6 757 36 927
rect 142 915 163 927
rect 216 915 237 927
rect 332 915 353 927
rect 75 826 106 915
rect 106 814 127 826
rect 180 814 201 826
rect 294 814 315 826
rect 370 814 391 826
rect 106 802 201 814
rect 255 793 391 814
rect 66 769 152 790
rect 185 769 275 781
rect 66 757 87 769
rect 185 757 201 769
rect 254 757 275 769
rect 6 668 30 757
rect 6 656 51 668
rect 104 656 125 668
rect 275 668 346 757
rect 144 656 165 668
rect 216 656 237 668
rect 6 644 237 656
rect 0 575 268 587
rect 349 571 353 590
rect 0 546 230 558
rect 251 546 295 558
rect 314 546 398 558
rect 0 517 398 529
rect 0 488 398 500
rect 0 459 92 471
rect 113 459 398 471
rect 0 430 204 442
rect 225 430 398 442
rect 6 364 165 376
rect 6 352 51 364
rect 144 352 165 364
rect 6 303 30 352
rect 275 303 346 352
rect 6 184 36 303
rect 104 278 125 303
rect 104 257 156 278
rect 257 257 317 278
rect 294 245 317 257
rect 75 196 106 245
rect 216 184 237 196
rect 370 184 391 196
rect 6 159 391 184
rect 6 36 36 159
rect 216 147 237 159
rect 332 147 353 159
rect 68 60 89 98
rect 256 86 277 98
rect 151 74 277 86
rect 68 48 308 60
rect 0 15 16 36
rect 37 15 68 36
rect 89 15 144 36
rect 165 15 218 36
rect 239 15 292 36
rect 313 15 369 36
rect 390 15 398 36
rect 0 6 398 15
<< m2contact >>
rect 330 571 349 590
rect 295 541 314 560
<< metal2 >>
rect 297 560 311 1182
rect 330 590 344 1182
rect 297 0 311 541
rect 330 0 344 571
<< labels >>
rlabel metal1 0 6 0 36 3 GND!
rlabel metal2 330 0 344 0 1 nQ
rlabel metal2 297 0 311 0 1 Q
rlabel metal1 398 6 398 36 7 GND!
rlabel metal1 0 459 0 471 1 Clock
rlabel metal1 0 430 0 442 1 nReset
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 546 0 558 1 Q
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 398 517 398 529 7 ScanReturn
rlabel metal1 398 546 398 558 7 Q
rlabel metal1 398 488 398 500 7 Test
rlabel metal1 398 459 398 471 7 Clock
rlabel metal1 398 430 398 442 7 nReset
rlabel metal1 0 575 0 587 1 nD
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel metal2 330 1182 344 1182 5 nQ
rlabel metal2 297 1182 311 1182 5 Q
rlabel metal1 398 1146 398 1176 7 Vdd!
<< end >>
