magic
tech tsmc180
timestamp 1733140770
<< nwell >>
rect 0 637 252 1176
<< polysilicon >>
rect 31 1119 40 1131
rect 69 1119 78 1131
rect 31 994 40 1030
rect 69 994 78 1030
rect 105 994 114 1131
rect 141 994 150 1131
rect 179 1119 188 1131
rect 224 1087 233 1131
rect 31 829 40 905
rect 31 198 40 802
rect 69 198 78 905
rect 105 869 114 905
rect 105 198 114 842
rect 141 828 150 905
rect 179 893 188 1030
rect 141 198 150 801
rect 179 255 188 872
rect 224 856 233 1066
rect 31 112 40 149
rect 69 112 78 149
rect 31 44 40 63
rect 69 44 78 63
rect 105 44 114 149
rect 141 44 150 149
rect 179 112 188 234
rect 224 101 233 829
rect 179 44 188 63
rect 224 44 233 80
<< ndiffusion >>
rect 28 149 31 198
rect 40 149 44 198
rect 65 149 69 198
rect 78 149 105 198
rect 114 149 117 198
rect 138 149 141 198
rect 150 149 153 198
rect 28 63 31 112
rect 40 63 43 112
rect 176 63 179 112
rect 188 63 191 112
<< pdiffusion >>
rect 28 1030 31 1119
rect 40 1030 43 1119
rect 176 1030 179 1119
rect 188 1030 191 1119
rect 28 905 31 994
rect 40 905 43 994
rect 64 905 69 994
rect 78 905 81 994
rect 102 905 105 994
rect 114 905 117 994
rect 138 905 141 994
rect 150 905 153 994
<< pohmic >>
rect 0 15 15 36
rect 36 15 101 36
rect 122 15 159 36
rect 180 15 205 36
rect 226 15 252 36
<< nohmic >>
rect 0 1146 20 1167
rect 41 1146 97 1167
rect 118 1146 162 1167
rect 183 1146 208 1167
rect 229 1146 252 1167
<< ntransistor >>
rect 31 149 40 198
rect 69 149 78 198
rect 105 149 114 198
rect 141 149 150 198
rect 31 63 40 112
rect 179 63 188 112
<< ptransistor >>
rect 31 1030 40 1119
rect 179 1030 188 1119
rect 31 905 40 994
rect 69 905 78 994
rect 105 905 114 994
rect 141 905 150 994
<< polycontact >>
rect 69 1030 90 1119
rect 224 1066 245 1087
rect 23 802 50 829
rect 91 842 118 869
rect 167 872 188 893
rect 128 801 155 828
rect 206 829 233 856
rect 167 234 188 255
rect 69 63 90 112
rect 224 80 245 101
<< ndiffcontact >>
rect 7 149 28 198
rect 44 149 65 198
rect 117 149 138 198
rect 153 149 174 198
rect 7 63 28 112
rect 43 63 64 112
rect 155 63 176 112
rect 191 63 212 112
<< pdiffcontact >>
rect 7 1030 28 1119
rect 43 1030 64 1119
rect 155 1030 176 1119
rect 191 1030 212 1119
rect 7 905 28 994
rect 43 905 64 994
rect 81 905 102 994
rect 117 905 138 994
rect 153 905 174 994
<< psubstratetap >>
rect 15 15 36 36
rect 101 15 122 36
rect 159 15 180 36
rect 205 15 226 36
<< nsubstratetap >>
rect 20 1146 41 1167
rect 97 1146 118 1167
rect 162 1146 183 1167
rect 208 1146 229 1167
<< metal1 >>
rect 0 1167 252 1176
rect 0 1146 20 1167
rect 41 1146 97 1167
rect 118 1146 162 1167
rect 183 1146 208 1167
rect 229 1146 252 1167
rect 7 1119 28 1146
rect 153 1119 174 1146
rect 64 1030 69 1119
rect 153 1030 155 1119
rect 212 1072 224 1084
rect 7 994 28 1030
rect 43 1006 138 1018
rect 43 994 64 1006
rect 117 994 138 1006
rect 153 994 174 1030
rect 86 893 98 905
rect 86 881 167 893
rect 0 546 252 558
rect 0 517 252 529
rect 0 488 252 500
rect 0 459 252 471
rect 0 430 252 442
rect 48 234 167 246
rect 48 198 60 234
rect 87 210 174 222
rect 7 137 28 149
rect 87 137 99 210
rect 153 198 174 210
rect 7 125 99 137
rect 64 63 69 112
rect 7 36 28 63
rect 117 36 138 149
rect 212 84 224 96
rect 155 36 176 63
rect 0 15 15 36
rect 36 15 101 36
rect 122 15 159 36
rect 180 15 205 36
rect 226 15 252 36
rect 0 6 252 15
<< m2contact >>
rect 91 842 118 869
rect 198 829 206 856
rect 206 829 225 856
rect 23 802 50 829
rect 128 801 155 828
<< metal2 >>
rect 33 829 47 1182
rect 99 869 113 1182
rect 33 0 47 802
rect 99 0 113 842
rect 132 828 146 1182
rect 198 856 212 1182
rect 132 0 146 801
rect 198 0 212 829
<< labels >>
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel metal1 0 546 0 558 3 SDI
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 430 0 442 3 nReset
rlabel metal1 0 6 0 36 3 GND!
rlabel metal1 252 1146 252 1176 7 Vdd!
rlabel metal1 252 6 252 36 7 GND!
rlabel metal2 33 1182 47 1182 5 S
rlabel metal2 33 0 47 0 1 S
rlabel metal2 99 0 113 0 1 I0
rlabel metal2 132 0 146 0 1 I1
rlabel metal2 198 0 212 0 1 Y
rlabel metal2 99 1182 113 1182 5 I0
rlabel metal2 132 1182 146 1182 5 I1
rlabel metal2 198 1182 212 1182 5 Y
rlabel metal1 252 546 252 558 7 SDI
rlabel metal1 252 517 252 529 7 ScanReturn
rlabel metal1 252 488 252 500 7 Test
rlabel metal1 252 459 252 471 7 Clock
rlabel metal1 252 430 252 442 7 nReset
<< end >>
