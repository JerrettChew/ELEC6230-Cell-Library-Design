magic
tech tsmc180
timestamp 1733141744
<< nwell >>
rect 454 637 2520 1176
<< polysilicon >>
rect 486 1119 495 1130
rect 601 1119 610 1130
rect 716 1119 725 1130
rect 831 1119 840 1130
rect 878 1119 887 1130
rect 979 1119 988 1130
rect 1027 1119 1036 1130
rect 1063 1119 1072 1130
rect 1112 1119 1121 1130
rect 1148 1119 1157 1130
rect 1262 1119 1271 1130
rect 1376 1119 1385 1130
rect 1491 1119 1500 1130
rect 1538 1119 1547 1130
rect 1639 1119 1648 1130
rect 1687 1119 1696 1130
rect 1723 1119 1732 1130
rect 1771 1119 1780 1130
rect 1807 1119 1816 1130
rect 1921 1119 1930 1130
rect 2036 1119 2045 1130
rect 2151 1119 2160 1130
rect 2198 1119 2207 1130
rect 2299 1119 2308 1130
rect 2347 1119 2356 1130
rect 2383 1119 2392 1130
rect 2431 1119 2440 1130
rect 2467 1119 2476 1130
rect 486 534 495 1030
rect 486 112 495 513
rect 601 505 610 1018
rect 716 505 725 846
rect 831 505 840 750
rect 601 100 610 484
rect 716 163 725 484
rect 831 231 840 484
rect 878 231 887 750
rect 979 505 988 716
rect 831 222 887 231
rect 831 198 840 222
rect 878 198 887 222
rect 979 231 988 484
rect 1027 231 1036 716
rect 1063 231 1072 716
rect 1112 231 1121 716
rect 1148 231 1157 716
rect 1262 476 1271 1018
rect 1376 476 1385 846
rect 1491 476 1500 750
rect 979 222 1157 231
rect 979 212 988 222
rect 1027 212 1036 222
rect 1063 212 1072 222
rect 1112 212 1121 222
rect 1148 212 1157 222
rect 1262 100 1271 455
rect 1376 163 1385 455
rect 1491 231 1500 455
rect 1538 231 1547 750
rect 1639 476 1648 716
rect 1491 222 1547 231
rect 1491 198 1500 222
rect 1538 198 1547 222
rect 1639 231 1648 455
rect 1687 231 1696 716
rect 1723 231 1732 716
rect 1771 231 1780 716
rect 1807 231 1816 716
rect 1921 447 1930 1018
rect 2036 447 2045 846
rect 2151 447 2160 750
rect 1639 222 1816 231
rect 1639 212 1648 222
rect 1687 212 1696 222
rect 1723 212 1732 222
rect 1771 212 1780 222
rect 1807 212 1816 222
rect 1921 100 1930 426
rect 2036 163 2045 426
rect 2151 231 2160 426
rect 2198 231 2207 750
rect 2299 447 2308 716
rect 2151 222 2207 231
rect 2151 198 2160 222
rect 2198 198 2207 222
rect 2299 231 2308 426
rect 2347 231 2356 716
rect 2383 231 2392 716
rect 2431 231 2440 716
rect 2467 231 2476 716
rect 2299 222 2476 231
rect 2299 212 2308 222
rect 2347 212 2356 222
rect 2383 212 2392 222
rect 2431 212 2440 222
rect 2467 212 2476 222
rect 486 52 495 63
rect 601 52 610 63
rect 716 52 725 63
rect 831 52 840 63
rect 878 52 887 63
rect 979 52 988 63
rect 1027 52 1036 63
rect 1063 52 1072 63
rect 1112 52 1121 63
rect 1148 52 1157 63
rect 1262 52 1271 63
rect 1376 52 1385 63
rect 1491 52 1500 63
rect 1538 52 1547 63
rect 1639 52 1648 63
rect 1687 52 1696 63
rect 1723 52 1732 63
rect 1771 52 1780 63
rect 1807 52 1816 63
rect 1921 52 1930 63
rect 2036 52 2045 63
rect 2151 52 2160 63
rect 2198 52 2207 63
rect 2299 52 2308 63
rect 2347 52 2356 63
rect 2383 52 2392 63
rect 2431 52 2440 63
rect 2467 52 2476 63
<< ndiffusion >>
rect 483 63 486 112
rect 495 63 498 112
rect 598 63 601 100
rect 610 63 613 100
rect 713 63 716 163
rect 725 63 728 163
rect 828 63 831 198
rect 840 63 843 198
rect 864 63 878 198
rect 887 63 890 198
rect 976 63 979 212
rect 988 63 991 212
rect 1012 63 1027 212
rect 1036 63 1039 212
rect 1060 63 1063 212
rect 1072 63 1075 212
rect 1096 63 1112 212
rect 1121 63 1124 212
rect 1145 63 1148 212
rect 1157 63 1160 212
rect 1259 63 1262 100
rect 1271 63 1274 100
rect 1373 63 1376 163
rect 1385 63 1388 163
rect 1488 63 1491 198
rect 1500 63 1503 198
rect 1524 63 1538 198
rect 1547 63 1550 198
rect 1636 63 1639 212
rect 1648 63 1651 212
rect 1672 63 1687 212
rect 1696 63 1699 212
rect 1720 63 1723 212
rect 1732 63 1735 212
rect 1756 63 1771 212
rect 1780 63 1783 212
rect 1804 63 1807 212
rect 1816 63 1819 212
rect 1918 63 1921 100
rect 1930 63 1933 100
rect 2033 63 2036 163
rect 2045 63 2048 163
rect 2148 63 2151 198
rect 2160 63 2163 198
rect 2184 63 2198 198
rect 2207 63 2210 198
rect 2296 63 2299 212
rect 2308 63 2311 212
rect 2332 63 2347 212
rect 2356 63 2359 212
rect 2380 63 2383 212
rect 2392 63 2395 212
rect 2416 63 2431 212
rect 2440 63 2443 212
rect 2464 63 2467 212
rect 2476 63 2479 212
<< pdiffusion >>
rect 483 1030 486 1119
rect 495 1030 498 1119
rect 598 1018 601 1119
rect 610 1018 613 1119
rect 713 846 716 1119
rect 725 846 728 1119
rect 828 750 831 1119
rect 840 750 843 1119
rect 864 750 878 1119
rect 887 750 890 1119
rect 976 716 979 1119
rect 988 716 991 1119
rect 1012 716 1027 1119
rect 1036 716 1039 1119
rect 1060 716 1063 1119
rect 1072 716 1075 1119
rect 1096 716 1112 1119
rect 1121 716 1124 1119
rect 1145 716 1148 1119
rect 1157 716 1160 1119
rect 1259 1018 1262 1119
rect 1271 1018 1274 1119
rect 1373 846 1376 1119
rect 1385 846 1388 1119
rect 1488 750 1491 1119
rect 1500 750 1503 1119
rect 1524 750 1538 1119
rect 1547 750 1550 1119
rect 1636 716 1639 1119
rect 1648 716 1651 1119
rect 1672 716 1687 1119
rect 1696 716 1699 1119
rect 1720 716 1723 1119
rect 1732 716 1735 1119
rect 1756 716 1771 1119
rect 1780 716 1783 1119
rect 1804 716 1807 1119
rect 1816 716 1819 1119
rect 1918 1018 1921 1119
rect 1930 1018 1933 1119
rect 2033 846 2036 1119
rect 2045 846 2048 1119
rect 2148 750 2151 1119
rect 2160 750 2163 1119
rect 2184 750 2198 1119
rect 2207 750 2210 1119
rect 2296 716 2299 1119
rect 2308 716 2311 1119
rect 2332 716 2347 1119
rect 2356 716 2359 1119
rect 2380 716 2383 1119
rect 2392 716 2395 1119
rect 2416 716 2431 1119
rect 2440 716 2443 1119
rect 2464 716 2467 1119
rect 2476 716 2479 1119
<< pohmic >>
rect 0 15 330 36
rect 351 15 396 36
rect 417 15 462 36
rect 483 15 577 36
rect 598 15 692 36
rect 713 15 807 36
rect 828 15 890 36
rect 911 15 955 36
rect 976 15 1039 36
rect 1060 15 1238 36
rect 1259 15 1352 36
rect 1373 15 1467 36
rect 1488 15 1550 36
rect 1571 15 1615 36
rect 1636 15 1699 36
rect 1720 15 1897 36
rect 1918 15 2012 36
rect 2033 15 2127 36
rect 2148 15 2210 36
rect 2231 15 2275 36
rect 2296 15 2359 36
rect 2380 15 2520 36
<< nohmic >>
rect 0 1146 33 1167
rect 54 1146 132 1167
rect 153 1146 231 1167
rect 252 1146 330 1167
rect 351 1146 396 1167
rect 417 1146 462 1167
rect 483 1146 577 1167
rect 598 1146 692 1167
rect 713 1146 807 1167
rect 828 1146 890 1167
rect 912 1146 955 1167
rect 976 1146 1039 1167
rect 1060 1146 1124 1167
rect 1145 1146 1238 1167
rect 1259 1146 1352 1167
rect 1373 1146 1467 1167
rect 1488 1146 1550 1167
rect 1572 1146 1615 1167
rect 1636 1146 1699 1167
rect 1720 1146 1783 1167
rect 1804 1146 1897 1167
rect 1918 1146 2012 1167
rect 2033 1146 2127 1167
rect 2148 1146 2210 1167
rect 2232 1146 2275 1167
rect 2296 1146 2359 1167
rect 2380 1146 2443 1167
rect 2464 1146 2520 1167
<< ntransistor >>
rect 486 63 495 112
rect 601 63 610 100
rect 716 63 725 163
rect 831 63 840 198
rect 878 63 887 198
rect 979 63 988 212
rect 1027 63 1036 212
rect 1063 63 1072 212
rect 1112 63 1121 212
rect 1148 63 1157 212
rect 1262 63 1271 100
rect 1376 63 1385 163
rect 1491 63 1500 198
rect 1538 63 1547 198
rect 1639 63 1648 212
rect 1687 63 1696 212
rect 1723 63 1732 212
rect 1771 63 1780 212
rect 1807 63 1816 212
rect 1921 63 1930 100
rect 2036 63 2045 163
rect 2151 63 2160 198
rect 2198 63 2207 198
rect 2299 63 2308 212
rect 2347 63 2356 212
rect 2383 63 2392 212
rect 2431 63 2440 212
rect 2467 63 2476 212
<< ptransistor >>
rect 486 1030 495 1119
rect 601 1018 610 1119
rect 716 846 725 1119
rect 831 750 840 1119
rect 878 750 887 1119
rect 979 716 988 1119
rect 1027 716 1036 1119
rect 1063 716 1072 1119
rect 1112 716 1121 1119
rect 1148 716 1157 1119
rect 1262 1018 1271 1119
rect 1376 846 1385 1119
rect 1491 750 1500 1119
rect 1538 750 1547 1119
rect 1639 716 1648 1119
rect 1687 716 1696 1119
rect 1723 716 1732 1119
rect 1771 716 1780 1119
rect 1807 716 1816 1119
rect 1921 1018 1930 1119
rect 2036 846 2045 1119
rect 2151 750 2160 1119
rect 2198 750 2207 1119
rect 2299 716 2308 1119
rect 2347 716 2356 1119
rect 2383 716 2392 1119
rect 2431 716 2440 1119
rect 2467 716 2476 1119
<< polycontact >>
rect 486 513 507 534
rect 589 484 610 505
rect 704 484 725 505
rect 819 484 840 505
rect 967 484 988 505
rect 1250 455 1271 476
rect 1364 455 1385 476
rect 1479 455 1500 476
rect 1627 455 1648 476
rect 1909 426 1930 447
rect 2024 426 2045 447
rect 2139 426 2160 447
rect 2287 426 2308 447
<< ndiffcontact >>
rect 462 63 483 112
rect 498 63 519 112
rect 577 63 598 100
rect 613 63 634 100
rect 692 63 713 163
rect 728 63 749 163
rect 807 63 828 198
rect 843 63 864 198
rect 890 63 911 198
rect 955 63 976 212
rect 991 63 1012 212
rect 1039 63 1060 212
rect 1075 63 1096 212
rect 1124 63 1145 212
rect 1160 63 1181 212
rect 1238 63 1259 100
rect 1274 63 1295 100
rect 1352 63 1373 163
rect 1388 63 1409 163
rect 1467 63 1488 198
rect 1503 63 1524 198
rect 1550 63 1571 198
rect 1615 63 1636 212
rect 1651 63 1672 212
rect 1699 63 1720 212
rect 1735 63 1756 212
rect 1783 63 1804 212
rect 1819 63 1840 212
rect 1897 63 1918 100
rect 1933 63 1954 100
rect 2012 63 2033 163
rect 2048 63 2069 163
rect 2127 63 2148 198
rect 2163 63 2184 198
rect 2210 63 2231 198
rect 2275 63 2296 212
rect 2311 63 2332 212
rect 2359 63 2380 212
rect 2395 63 2416 212
rect 2443 63 2464 212
rect 2479 63 2500 212
<< pdiffcontact >>
rect 462 1030 483 1119
rect 498 1030 519 1119
rect 577 1018 598 1119
rect 613 1018 634 1119
rect 692 846 713 1119
rect 728 846 749 1119
rect 807 750 828 1119
rect 843 750 864 1119
rect 890 750 911 1119
rect 955 716 976 1119
rect 991 716 1012 1119
rect 1039 716 1060 1119
rect 1075 716 1096 1119
rect 1124 716 1145 1119
rect 1160 716 1181 1119
rect 1238 1018 1259 1119
rect 1274 1018 1295 1119
rect 1352 846 1373 1119
rect 1388 846 1409 1119
rect 1467 750 1488 1119
rect 1503 750 1524 1119
rect 1550 750 1571 1119
rect 1615 716 1636 1119
rect 1651 716 1672 1119
rect 1699 716 1720 1119
rect 1735 716 1756 1119
rect 1783 716 1804 1119
rect 1819 716 1840 1119
rect 1897 1018 1918 1119
rect 1933 1018 1954 1119
rect 2012 846 2033 1119
rect 2048 846 2069 1119
rect 2127 750 2148 1119
rect 2163 750 2184 1119
rect 2210 750 2231 1119
rect 2275 716 2296 1119
rect 2311 716 2332 1119
rect 2359 716 2380 1119
rect 2395 716 2416 1119
rect 2443 716 2464 1119
rect 2479 716 2500 1119
<< psubstratetap >>
rect 330 15 351 36
rect 396 15 417 36
rect 462 15 483 36
rect 577 15 598 36
rect 692 15 713 36
rect 807 15 828 36
rect 890 15 911 36
rect 955 15 976 36
rect 1039 15 1060 36
rect 1238 15 1259 36
rect 1352 15 1373 36
rect 1467 15 1488 36
rect 1550 15 1571 36
rect 1615 15 1636 36
rect 1699 15 1720 36
rect 1897 15 1918 36
rect 2012 15 2033 36
rect 2127 15 2148 36
rect 2210 15 2231 36
rect 2275 15 2296 36
rect 2359 15 2380 36
<< nsubstratetap >>
rect 33 1146 54 1167
rect 132 1146 153 1167
rect 231 1146 252 1167
rect 330 1146 351 1167
rect 396 1146 417 1167
rect 462 1146 483 1167
rect 577 1146 598 1167
rect 692 1146 713 1167
rect 807 1146 828 1167
rect 890 1146 912 1167
rect 955 1146 976 1167
rect 1039 1146 1060 1167
rect 1124 1146 1145 1167
rect 1238 1146 1259 1167
rect 1352 1146 1373 1167
rect 1467 1146 1488 1167
rect 1550 1146 1572 1167
rect 1615 1146 1636 1167
rect 1699 1146 1720 1167
rect 1783 1146 1804 1167
rect 1897 1146 1918 1167
rect 2012 1146 2033 1167
rect 2127 1146 2148 1167
rect 2210 1146 2232 1167
rect 2275 1146 2296 1167
rect 2359 1146 2380 1167
rect 2443 1146 2464 1167
<< metal1 >>
rect 300 1167 2520 1176
rect 300 1146 330 1167
rect 351 1146 396 1167
rect 417 1146 462 1167
rect 483 1146 577 1167
rect 598 1146 692 1167
rect 713 1146 807 1167
rect 828 1146 890 1167
rect 912 1146 955 1167
rect 976 1146 1039 1167
rect 1060 1146 1124 1167
rect 1145 1146 1238 1167
rect 1259 1146 1352 1167
rect 1373 1146 1467 1167
rect 1488 1146 1550 1167
rect 1572 1146 1615 1167
rect 1636 1146 1699 1167
rect 1720 1146 1783 1167
rect 1804 1146 1897 1167
rect 1918 1146 2012 1167
rect 2033 1146 2127 1167
rect 2148 1146 2210 1167
rect 2232 1146 2275 1167
rect 2296 1146 2359 1167
rect 2380 1146 2443 1167
rect 2464 1146 2520 1167
rect 462 1119 483 1146
rect 577 1119 598 1146
rect 692 1119 713 1146
rect 807 1119 828 1146
rect 890 1119 911 1146
rect 349 969 512 981
rect 955 1119 976 1146
rect 1039 1119 1060 1146
rect 1124 1119 1145 1146
rect 1238 1119 1259 1146
rect 1352 1119 1373 1146
rect 1467 1119 1488 1146
rect 1550 1119 1571 1146
rect 1615 1119 1636 1146
rect 1699 1119 1720 1146
rect 1783 1119 1804 1146
rect 1897 1119 1918 1146
rect 2012 1119 2033 1146
rect 2127 1119 2148 1146
rect 2210 1119 2231 1146
rect 2275 1119 2296 1146
rect 2359 1119 2380 1146
rect 2443 1119 2464 1146
rect 347 546 2520 558
rect 507 517 2520 529
rect 382 488 589 500
rect 648 488 704 500
rect 763 488 819 500
rect 877 488 967 500
rect 1194 488 2520 500
rect 415 459 1250 471
rect 1309 459 1364 471
rect 1423 459 1479 471
rect 1537 459 1627 471
rect 1853 459 2520 471
rect 448 430 1909 442
rect 1968 430 2024 442
rect 2083 430 2139 442
rect 2197 430 2287 442
rect 2513 430 2520 442
rect 462 36 483 63
rect 577 36 598 63
rect 692 36 713 63
rect 807 36 828 63
rect 890 36 911 63
rect 955 36 976 63
rect 1039 36 1060 63
rect 1124 36 1145 63
rect 1238 36 1259 63
rect 1352 36 1373 63
rect 1467 36 1488 63
rect 1550 36 1571 63
rect 1615 36 1636 63
rect 1699 36 1720 63
rect 1783 36 1804 63
rect 1897 36 1918 63
rect 2012 36 2033 63
rect 2127 36 2148 63
rect 2210 36 2231 63
rect 2275 36 2296 63
rect 2359 36 2380 63
rect 2443 36 2464 63
rect 0 15 330 36
rect 351 15 396 36
rect 417 15 462 36
rect 483 15 577 36
rect 598 15 692 36
rect 713 15 807 36
rect 828 15 890 36
rect 911 15 955 36
rect 976 15 1039 36
rect 1060 15 1238 36
rect 1259 15 1352 36
rect 1373 15 1467 36
rect 1488 15 1550 36
rect 1571 15 1615 36
rect 1636 15 1699 36
rect 1720 15 1897 36
rect 1918 15 2012 36
rect 2033 15 2127 36
rect 2148 15 2210 36
rect 2231 15 2275 36
rect 2296 15 2359 36
rect 2380 15 2520 36
rect 0 6 2520 15
<< m2contact >>
rect 0 1167 300 1176
rect 0 1146 33 1167
rect 33 1146 54 1167
rect 54 1146 132 1167
rect 132 1146 153 1167
rect 153 1146 231 1167
rect 231 1146 252 1167
rect 252 1146 300 1167
rect 511 1030 519 1119
rect 519 1030 532 1119
rect 626 1018 634 1119
rect 634 1018 647 1119
rect 330 967 349 986
rect 512 965 533 986
rect 741 846 749 1119
rect 749 846 762 1119
rect 853 750 864 1119
rect 864 750 874 1119
rect 1002 716 1012 1119
rect 1012 716 1023 1119
rect 1086 716 1096 1119
rect 1096 716 1107 1119
rect 1171 716 1181 1119
rect 1181 716 1192 1119
rect 1287 1018 1295 1119
rect 1295 1018 1308 1119
rect 1401 846 1409 1119
rect 1409 846 1422 1119
rect 1513 750 1524 1119
rect 1524 750 1534 1119
rect 1662 716 1672 1119
rect 1672 716 1683 1119
rect 1746 716 1756 1119
rect 1756 716 1767 1119
rect 1830 716 1840 1119
rect 1840 716 1851 1119
rect 1946 1018 1954 1119
rect 1954 1018 1967 1119
rect 2061 846 2069 1119
rect 2069 846 2082 1119
rect 2173 750 2184 1119
rect 2184 750 2194 1119
rect 2322 716 2332 1119
rect 2332 716 2343 1119
rect 2406 716 2416 1119
rect 2416 716 2427 1119
rect 2490 716 2500 1119
rect 2500 716 2511 1119
rect 328 543 347 562
rect 363 485 382 504
rect 627 484 648 505
rect 742 484 763 505
rect 856 483 877 504
rect 1173 483 1194 504
rect 396 456 415 475
rect 1288 455 1309 476
rect 1402 455 1423 476
rect 1516 455 1537 476
rect 1832 454 1853 475
rect 429 427 448 446
rect 1947 425 1968 446
rect 2062 425 2083 446
rect 2176 425 2197 446
rect 2492 425 2513 446
rect 511 63 519 112
rect 519 63 532 112
rect 626 63 634 100
rect 634 63 647 100
rect 741 63 749 163
rect 749 63 762 163
rect 853 63 864 198
rect 864 63 874 198
rect 1003 63 1012 212
rect 1012 63 1024 212
rect 1086 63 1096 212
rect 1096 63 1107 212
rect 1171 63 1181 212
rect 1181 63 1192 212
rect 1287 63 1295 100
rect 1295 63 1308 100
rect 1401 63 1409 163
rect 1409 63 1422 163
rect 1513 63 1524 198
rect 1524 63 1534 198
rect 1663 63 1672 212
rect 1672 63 1684 212
rect 1746 63 1756 212
rect 1756 63 1767 212
rect 1830 63 1840 212
rect 1840 63 1851 212
rect 1946 63 1954 100
rect 1954 63 1967 100
rect 2061 63 2069 163
rect 2069 63 2082 163
rect 2173 63 2184 198
rect 2184 63 2194 198
rect 2323 63 2332 212
rect 2332 63 2344 212
rect 2406 63 2416 212
rect 2416 63 2427 212
rect 2490 63 2500 212
rect 2500 63 2511 212
<< metal2 >>
rect 0 1176 300 1182
rect 0 0 300 1146
rect 330 986 344 1182
rect 330 0 344 543
rect 363 504 377 1182
rect 363 0 377 485
rect 396 475 410 1182
rect 396 0 410 456
rect 429 446 443 1182
rect 512 1119 533 1130
rect 627 1119 648 1130
rect 742 1119 763 1130
rect 856 1119 877 1130
rect 1005 1119 1026 1130
rect 1089 1119 1110 1130
rect 1173 1119 1194 1130
rect 1288 1119 1309 1130
rect 1402 1119 1423 1130
rect 1516 1119 1537 1130
rect 1665 1119 1686 1130
rect 1749 1119 1770 1130
rect 1832 1119 1853 1130
rect 1947 1119 1968 1130
rect 2062 1119 2083 1130
rect 2176 1119 2197 1130
rect 2325 1119 2346 1130
rect 2409 1119 2430 1130
rect 2492 1119 2513 1130
rect 532 1030 533 1119
rect 512 986 533 1030
rect 647 1018 648 1119
rect 429 0 443 427
rect 512 112 533 965
rect 532 63 533 112
rect 627 505 648 1018
rect 762 846 763 1119
rect 627 100 648 484
rect 742 505 763 846
rect 874 750 877 1119
rect 742 163 763 484
rect 856 504 877 750
rect 1023 716 1026 1119
rect 1107 716 1110 1119
rect 1192 716 1194 1119
rect 1308 1018 1309 1119
rect 856 198 877 483
rect 1005 264 1026 716
rect 1089 264 1110 716
rect 1173 504 1194 716
rect 1173 264 1194 483
rect 1005 243 1194 264
rect 1005 212 1026 243
rect 1089 212 1110 243
rect 1173 212 1194 243
rect 647 63 648 100
rect 762 63 763 163
rect 874 63 877 198
rect 1024 63 1026 212
rect 1107 63 1110 212
rect 1192 63 1194 212
rect 1288 476 1309 1018
rect 1422 846 1423 1119
rect 1288 100 1309 455
rect 1402 476 1423 846
rect 1534 750 1537 1119
rect 1402 163 1423 455
rect 1516 476 1537 750
rect 1683 716 1686 1119
rect 1767 716 1770 1119
rect 1851 716 1853 1119
rect 1967 1018 1968 1119
rect 1516 198 1537 455
rect 1665 264 1686 716
rect 1749 264 1770 716
rect 1832 475 1853 716
rect 1832 264 1853 454
rect 1665 243 1853 264
rect 1665 212 1686 243
rect 1749 212 1770 243
rect 1832 212 1853 243
rect 1308 63 1309 100
rect 1422 63 1423 163
rect 1534 63 1537 198
rect 1684 63 1686 212
rect 1767 63 1770 212
rect 1851 63 1853 212
rect 1947 446 1968 1018
rect 2082 846 2083 1119
rect 1947 100 1968 425
rect 2062 446 2083 846
rect 2194 750 2197 1119
rect 2062 163 2083 425
rect 2176 446 2197 750
rect 2343 716 2346 1119
rect 2427 716 2430 1119
rect 2511 716 2513 1119
rect 2176 198 2197 425
rect 2325 264 2346 716
rect 2409 264 2430 716
rect 2492 446 2513 716
rect 2492 264 2513 425
rect 2325 243 2513 264
rect 2325 212 2346 243
rect 2409 212 2430 243
rect 2492 212 2513 243
rect 1967 63 1968 100
rect 2082 63 2083 163
rect 2194 63 2197 198
rect 2344 63 2346 212
rect 2427 63 2430 212
rect 2511 63 2513 212
rect 512 52 533 63
rect 627 52 648 63
rect 742 52 763 63
rect 856 52 877 63
rect 1005 52 1026 63
rect 1089 52 1110 63
rect 1173 52 1194 63
rect 1288 52 1309 63
rect 1402 52 1423 63
rect 1516 52 1537 63
rect 1665 52 1686 63
rect 1749 52 1770 63
rect 1832 52 1853 63
rect 1947 52 1968 63
rect 2062 52 2083 63
rect 2176 52 2197 63
rect 2325 52 2346 63
rect 2409 52 2430 63
rect 2492 52 2513 63
<< labels >>
rlabel metal2 0 0 300 0 1 Vdd!
rlabel metal2 0 1182 300 1182 5 Vdd!
rlabel metal2 363 1182 377 1182 5 Test
rlabel metal2 330 1182 344 1182 5 SDO
rlabel metal2 429 0 443 0 1 nReset
rlabel metal2 330 0 344 0 1 SDI
rlabel metal2 363 0 377 0 1 Test
rlabel metal2 396 0 410 0 1 Clock
rlabel metal1 2520 517 2520 529 7 nSDO
rlabel metal1 2520 430 2520 442 1 nResetOut
rlabel metal1 2520 459 2520 471 1 ClockOut
rlabel metal1 2520 488 2520 500 1 TestOut
rlabel metal1 2520 1146 2520 1176 1 Vdd!
rlabel metal1 2520 6 2520 36 7 GND!
rlabel metal2 396 1182 410 1182 5 Clock
rlabel metal2 429 1182 443 1182 5 nReset
rlabel metal1 2520 546 2520 558 7 SDI
rlabel metal1 0 6 0 36 1 GND!
<< end >>
