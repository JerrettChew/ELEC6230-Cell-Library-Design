magic
tech tsmc180
timestamp 1733141518
<< nwell >>
rect 0 637 789 1176
<< polysilicon >>
rect 31 994 40 1133
rect 142 1119 151 1133
rect 71 994 80 1030
rect 142 994 151 1030
rect 180 994 189 1133
rect 218 1119 227 1133
rect 218 994 227 1030
rect 289 994 298 1133
rect 325 994 334 1030
rect 373 994 382 1134
rect 445 915 454 1141
rect 483 1053 492 1141
rect 521 1110 530 1141
rect 521 1089 525 1110
rect 521 1053 530 1089
rect 559 1053 568 1141
rect 595 1053 604 1141
rect 31 591 40 905
rect 31 200 40 570
rect 71 200 80 905
rect 142 845 151 905
rect 180 845 189 905
rect 142 200 151 824
rect 180 200 189 824
rect 218 504 227 905
rect 289 563 298 905
rect 218 200 227 483
rect 289 200 298 542
rect 325 233 334 905
rect 373 869 382 905
rect 373 592 382 848
rect 445 757 454 826
rect 483 757 492 964
rect 521 915 530 964
rect 559 915 568 964
rect 595 915 604 964
rect 373 299 382 571
rect 445 352 454 668
rect 483 475 492 668
rect 483 352 492 454
rect 325 200 334 212
rect 31 44 40 151
rect 71 112 80 151
rect 142 112 151 151
rect 142 44 151 63
rect 180 44 189 151
rect 218 112 227 151
rect 218 44 227 63
rect 289 44 298 151
rect 325 44 334 151
rect 372 44 381 278
rect 445 245 454 303
rect 445 41 454 196
rect 483 147 492 303
rect 521 245 530 826
rect 559 790 568 826
rect 564 769 568 790
rect 559 757 568 769
rect 595 757 604 826
rect 633 814 642 1141
rect 671 1053 680 1141
rect 711 1134 720 1141
rect 711 1053 720 1113
rect 633 757 642 793
rect 559 352 568 668
rect 595 446 604 668
rect 633 562 642 668
rect 671 593 680 964
rect 711 915 720 964
rect 749 915 758 1141
rect 595 352 604 425
rect 633 352 642 541
rect 559 278 568 303
rect 559 245 568 257
rect 595 245 604 303
rect 633 278 642 303
rect 521 147 530 196
rect 559 147 568 196
rect 595 147 604 196
rect 483 41 492 98
rect 521 93 530 98
rect 521 41 530 72
rect 559 41 568 98
rect 595 41 604 98
rect 633 41 642 257
rect 671 147 680 572
rect 711 245 720 826
rect 749 757 758 826
rect 749 591 758 668
rect 749 352 758 570
rect 749 245 758 303
rect 711 147 720 196
rect 671 41 680 98
rect 711 69 720 98
rect 711 41 720 48
rect 749 41 758 196
<< ndiffusion >>
rect 442 303 445 352
rect 454 303 483 352
rect 492 303 495 352
rect 28 151 31 200
rect 40 151 71 200
rect 80 151 93 200
rect 114 151 142 200
rect 151 151 180 200
rect 189 151 192 200
rect 213 151 218 200
rect 227 151 289 200
rect 298 151 301 200
rect 322 151 325 200
rect 334 151 346 200
rect 139 63 142 112
rect 151 63 154 112
rect 215 63 218 112
rect 227 63 263 112
rect 556 303 559 352
rect 568 303 595 352
rect 604 303 633 352
rect 642 303 645 352
rect 518 196 521 245
rect 530 196 559 245
rect 568 196 595 245
rect 604 196 607 245
rect 480 98 483 147
rect 492 98 521 147
rect 530 98 559 147
rect 568 98 595 147
rect 604 98 607 147
rect 708 196 711 245
rect 720 196 749 245
rect 758 196 761 245
rect 668 98 671 147
rect 680 98 711 147
rect 720 98 723 147
<< pdiffusion >>
rect 139 1030 142 1119
rect 151 1030 154 1119
rect 215 1030 218 1119
rect 227 1030 263 1119
rect 28 905 31 994
rect 40 905 45 994
rect 66 905 71 994
rect 80 905 83 994
rect 139 905 142 994
rect 151 905 155 994
rect 176 905 180 994
rect 189 905 194 994
rect 215 905 218 994
rect 227 905 230 994
rect 251 905 289 994
rect 298 905 301 994
rect 322 905 325 994
rect 334 905 337 994
rect 480 964 483 1053
rect 492 964 495 1053
rect 516 964 521 1053
rect 530 964 533 1053
rect 554 964 559 1053
rect 568 964 571 1053
rect 592 964 595 1053
rect 604 964 607 1053
rect 518 826 521 915
rect 530 826 533 915
rect 554 826 559 915
rect 568 826 571 915
rect 592 826 595 915
rect 604 826 607 915
rect 442 668 445 757
rect 454 668 457 757
rect 478 668 483 757
rect 492 668 495 757
rect 668 964 671 1053
rect 680 964 683 1053
rect 704 964 711 1053
rect 720 964 723 1053
rect 556 668 559 757
rect 568 668 571 757
rect 592 668 595 757
rect 604 668 607 757
rect 628 668 633 757
rect 642 668 645 757
rect 706 826 711 915
rect 720 826 723 915
rect 744 826 749 915
rect 758 826 761 915
<< pohmic >>
rect 0 15 44 36
rect 65 15 99 36
rect 120 15 194 36
rect 215 15 253 36
rect 274 15 301 36
rect 322 15 344 36
rect 365 15 407 36
rect 428 15 459 36
rect 480 15 535 36
rect 556 15 609 36
rect 630 15 683 36
rect 704 15 760 36
rect 781 15 789 36
<< nohmic >>
rect 0 1146 49 1167
rect 70 1146 109 1167
rect 130 1146 185 1167
rect 206 1146 231 1167
rect 252 1146 304 1167
rect 325 1146 360 1167
rect 381 1146 414 1167
rect 435 1146 457 1167
rect 478 1146 535 1167
rect 556 1146 608 1167
rect 629 1146 687 1167
rect 708 1146 759 1167
rect 780 1146 789 1167
<< ntransistor >>
rect 445 303 454 352
rect 483 303 492 352
rect 31 151 40 200
rect 71 151 80 200
rect 142 151 151 200
rect 180 151 189 200
rect 218 151 227 200
rect 289 151 298 200
rect 325 151 334 200
rect 142 63 151 112
rect 218 63 227 112
rect 559 303 568 352
rect 595 303 604 352
rect 633 303 642 352
rect 521 196 530 245
rect 559 196 568 245
rect 595 196 604 245
rect 483 98 492 147
rect 521 98 530 147
rect 559 98 568 147
rect 595 98 604 147
rect 711 196 720 245
rect 749 196 758 245
rect 671 98 680 147
rect 711 98 720 147
<< ptransistor >>
rect 142 1030 151 1119
rect 218 1030 227 1119
rect 31 905 40 994
rect 71 905 80 994
rect 142 905 151 994
rect 180 905 189 994
rect 218 905 227 994
rect 289 905 298 994
rect 325 905 334 994
rect 483 964 492 1053
rect 521 964 530 1053
rect 559 964 568 1053
rect 595 964 604 1053
rect 521 826 530 915
rect 559 826 568 915
rect 595 826 604 915
rect 445 668 454 757
rect 483 668 492 757
rect 671 964 680 1053
rect 711 964 720 1053
rect 559 668 568 757
rect 595 668 604 757
rect 633 668 642 757
rect 711 826 720 915
rect 749 826 758 915
<< polycontact >>
rect 71 1030 92 1119
rect 313 1030 334 1119
rect 363 905 384 994
rect 525 1089 546 1110
rect 25 570 46 591
rect 132 824 153 845
rect 174 824 195 845
rect 277 542 298 563
rect 212 483 233 504
rect 361 848 382 869
rect 445 826 466 915
rect 361 571 382 592
rect 483 454 504 475
rect 361 278 382 299
rect 313 212 334 233
rect 71 63 92 112
rect 445 196 466 245
rect 543 769 564 790
rect 699 1113 720 1134
rect 625 793 646 814
rect 659 572 680 593
rect 621 541 642 562
rect 595 425 616 446
rect 547 257 568 278
rect 627 257 648 278
rect 521 72 542 93
rect 737 668 758 757
rect 744 570 765 591
rect 737 303 758 352
rect 699 48 720 69
<< ndiffcontact >>
rect 421 303 442 352
rect 495 303 516 352
rect 7 151 28 200
rect 93 151 114 200
rect 192 151 213 200
rect 301 151 322 200
rect 346 151 367 200
rect 118 63 139 112
rect 154 63 175 112
rect 194 63 215 112
rect 263 63 284 112
rect 535 303 556 352
rect 645 303 666 352
rect 497 196 518 245
rect 607 196 628 245
rect 459 98 480 147
rect 607 98 628 147
rect 685 196 708 245
rect 761 196 782 245
rect 647 98 668 147
rect 723 98 744 147
<< pdiffcontact >>
rect 118 1030 139 1119
rect 154 1030 175 1119
rect 194 1030 215 1119
rect 263 1030 284 1119
rect 7 905 28 994
rect 45 905 66 994
rect 83 905 104 994
rect 118 905 139 994
rect 155 905 176 994
rect 194 905 215 994
rect 230 905 251 994
rect 301 905 322 994
rect 337 905 358 994
rect 459 964 480 1053
rect 495 964 516 1053
rect 533 964 554 1053
rect 571 964 592 1053
rect 607 964 628 1053
rect 497 826 518 915
rect 533 826 554 915
rect 571 826 592 915
rect 607 826 628 915
rect 421 668 442 757
rect 457 668 478 757
rect 495 668 516 757
rect 647 964 668 1053
rect 683 964 704 1053
rect 723 964 744 1053
rect 535 668 556 757
rect 571 668 592 757
rect 607 668 628 757
rect 645 668 666 757
rect 685 826 706 915
rect 723 826 744 915
rect 761 826 782 915
<< psubstratetap >>
rect 44 15 65 36
rect 99 15 120 36
rect 194 15 215 36
rect 253 15 274 36
rect 301 15 322 36
rect 344 15 365 36
rect 407 15 428 36
rect 459 15 480 36
rect 535 15 556 36
rect 609 15 630 36
rect 683 15 704 36
rect 760 15 781 36
<< nsubstratetap >>
rect 49 1146 70 1167
rect 109 1146 130 1167
rect 185 1146 206 1167
rect 231 1146 252 1167
rect 304 1146 325 1167
rect 360 1146 381 1167
rect 414 1146 435 1167
rect 457 1146 478 1167
rect 535 1146 556 1167
rect 608 1146 629 1167
rect 687 1146 708 1167
rect 759 1146 780 1167
<< metal1 >>
rect 0 1167 789 1176
rect 0 1146 49 1167
rect 70 1146 109 1167
rect 130 1146 185 1167
rect 206 1146 231 1167
rect 252 1146 304 1167
rect 325 1146 360 1167
rect 381 1146 414 1167
rect 435 1146 457 1167
rect 478 1146 535 1167
rect 556 1146 608 1167
rect 629 1146 687 1167
rect 708 1146 759 1167
rect 780 1146 789 1167
rect 154 1119 175 1146
rect 92 1030 118 1119
rect 194 1119 215 1146
rect 7 1006 104 1018
rect 7 994 28 1006
rect 83 994 104 1006
rect 45 869 66 905
rect 118 1006 215 1018
rect 118 994 139 1006
rect 194 994 215 1006
rect 230 994 251 1146
rect 284 1030 313 1119
rect 358 905 363 994
rect 397 952 427 1146
rect 495 1122 699 1134
rect 495 1077 513 1122
rect 546 1089 704 1101
rect 495 1065 592 1077
rect 495 1053 516 1065
rect 571 1053 592 1065
rect 683 1053 704 1089
rect 459 952 480 964
rect 533 952 554 964
rect 607 952 628 964
rect 647 952 668 964
rect 723 952 744 964
rect 397 927 744 952
rect 83 893 104 905
rect 155 893 175 905
rect 83 881 175 893
rect 194 893 215 905
rect 301 893 322 905
rect 194 881 322 893
rect 45 857 361 869
rect 397 757 427 927
rect 533 915 554 927
rect 607 915 628 927
rect 723 915 744 927
rect 466 826 497 915
rect 497 814 518 826
rect 571 814 592 826
rect 685 814 706 826
rect 761 814 782 826
rect 497 802 592 814
rect 646 793 782 814
rect 457 769 543 790
rect 576 769 666 781
rect 457 757 478 769
rect 576 757 592 769
rect 645 757 666 769
rect 397 668 421 757
rect 397 656 442 668
rect 495 656 516 668
rect 666 668 737 757
rect 535 656 556 668
rect 607 656 628 668
rect 397 644 628 656
rect 46 575 322 587
rect 0 546 277 558
rect 310 558 322 575
rect 382 575 659 587
rect 742 571 744 590
rect 310 546 621 558
rect 642 546 690 558
rect 709 546 789 558
rect 0 517 789 529
rect 0 488 212 500
rect 233 488 789 500
rect 0 459 483 471
rect 504 459 789 471
rect 0 430 595 442
rect 616 430 789 442
rect 397 364 556 376
rect 397 352 442 364
rect 535 352 556 364
rect 397 303 421 352
rect 666 303 737 352
rect 7 278 361 290
rect 7 200 28 278
rect 93 245 367 266
rect 93 200 114 245
rect 263 214 313 231
rect 7 139 28 151
rect 192 139 213 151
rect 7 124 213 139
rect 263 112 284 214
rect 346 200 367 245
rect 92 63 118 112
rect 154 36 175 63
rect 397 184 427 303
rect 495 278 516 303
rect 495 257 547 278
rect 648 257 708 278
rect 685 245 708 257
rect 466 196 497 245
rect 607 184 628 196
rect 761 184 782 196
rect 397 159 782 184
rect 194 36 215 63
rect 301 36 322 151
rect 397 36 427 159
rect 607 147 628 159
rect 723 147 744 159
rect 459 60 480 98
rect 647 86 668 98
rect 542 74 668 86
rect 459 48 699 60
rect 0 15 44 36
rect 65 15 99 36
rect 120 15 194 36
rect 215 15 253 36
rect 274 15 301 36
rect 322 15 344 36
rect 365 15 407 36
rect 428 15 459 36
rect 480 15 535 36
rect 556 15 609 36
rect 630 15 683 36
rect 704 15 760 36
rect 781 15 789 36
rect 0 6 789 15
<< m2contact >>
rect 124 824 132 845
rect 132 824 143 845
rect 165 824 174 845
rect 174 824 184 845
rect 723 571 742 590
rect 690 541 709 560
<< metal2 >>
rect 132 845 146 1182
rect 143 824 146 845
rect 132 0 146 824
rect 165 845 179 1182
rect 165 0 179 824
rect 693 560 707 1182
rect 726 590 740 1182
rect 693 0 707 541
rect 726 0 740 571
<< labels >>
rlabel metal2 132 1182 146 1182 5 Load
rlabel metal2 165 1182 179 1182 5 D
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 0 546 0 558 3 SDI
rlabel metal1 0 430 0 442 3 nReset
rlabel metal2 165 0 179 0 1 D
rlabel metal2 132 0 146 0 1 Load
rlabel metal1 0 6 0 36 3 GND!
rlabel metal1 789 6 789 36 7 GND!
rlabel metal1 789 517 789 529 7 ScanReturn
rlabel metal1 789 546 789 558 7 Q
rlabel metal1 789 488 789 500 7 Test
rlabel metal1 789 459 789 471 7 Clock
rlabel metal1 789 430 789 442 7 nReset
rlabel metal2 726 0 740 0 1 nQ
rlabel metal2 726 1182 740 1182 5 nQ
rlabel metal2 693 1182 707 1182 5 Q
rlabel metal2 693 0 707 0 1 Q
rlabel metal1 789 1146 789 1176 7 Vdd!
<< end >>
