magic
tech tsmc180
timestamp 1733140494
<< nwell >>
rect 0 637 291 1176
<< polysilicon >>
rect 66 1110 75 1126
rect 102 1110 111 1126
rect 173 1110 182 1121
rect 220 1110 229 1121
rect 66 948 75 1021
rect 102 948 111 1021
rect 173 1007 182 1021
rect 173 948 182 986
rect 66 846 75 859
rect 66 255 75 825
rect 102 823 111 859
rect 102 255 111 800
rect 173 255 182 859
rect 220 847 229 1021
rect 220 288 229 826
rect 66 122 75 206
rect 102 122 111 206
rect 173 179 182 206
rect 173 122 182 158
rect 220 122 229 267
rect 66 62 75 73
rect 102 62 111 73
rect 173 62 182 73
rect 220 62 229 73
<< ndiffusion >>
rect 63 206 66 255
rect 75 206 78 255
rect 99 206 102 255
rect 111 206 114 255
rect 135 206 173 255
rect 182 206 194 255
rect 63 73 66 122
rect 75 73 102 122
rect 111 73 114 122
rect 170 73 173 122
rect 182 73 194 122
rect 215 73 220 122
rect 229 73 232 122
<< pdiffusion >>
rect 63 1021 66 1110
rect 75 1021 78 1110
rect 99 1021 102 1110
rect 111 1021 114 1110
rect 170 1021 173 1110
rect 182 1021 194 1110
rect 215 1021 220 1110
rect 229 1021 232 1110
rect 63 859 66 948
rect 75 859 102 948
rect 111 859 114 948
rect 135 859 173 948
rect 182 859 194 948
<< pohmic >>
rect 0 15 2 36
rect 23 15 33 36
rect 54 15 66 36
rect 87 15 99 36
rect 120 15 132 36
rect 153 15 165 36
rect 186 15 198 36
rect 219 15 231 36
rect 252 15 264 36
rect 285 15 291 36
<< nohmic >>
rect 0 1146 2 1167
rect 23 1146 33 1167
rect 54 1146 66 1167
rect 87 1146 99 1167
rect 120 1146 132 1167
rect 153 1146 165 1167
rect 186 1146 198 1167
rect 219 1146 231 1167
rect 252 1146 264 1167
rect 285 1146 291 1167
<< ntransistor >>
rect 66 206 75 255
rect 102 206 111 255
rect 173 206 182 255
rect 66 73 75 122
rect 102 73 111 122
rect 173 73 182 122
rect 220 73 229 122
<< ptransistor >>
rect 66 1021 75 1110
rect 102 1021 111 1110
rect 173 1021 182 1110
rect 220 1021 229 1110
rect 66 859 75 948
rect 102 859 111 948
rect 173 859 182 948
<< polycontact >>
rect 161 986 182 1007
rect 60 825 81 846
rect 96 800 119 823
rect 211 826 232 847
rect 214 267 235 288
rect 161 158 182 179
<< ndiffcontact >>
rect 42 206 63 255
rect 78 206 99 255
rect 114 206 135 255
rect 194 206 215 255
rect 42 73 63 122
rect 114 73 135 122
rect 149 73 170 122
rect 194 73 215 122
rect 232 73 253 122
<< pdiffcontact >>
rect 42 1021 63 1110
rect 78 1021 99 1110
rect 114 1021 135 1110
rect 149 1021 170 1110
rect 194 1021 215 1110
rect 232 1021 253 1110
rect 42 859 63 948
rect 114 859 135 948
rect 194 859 215 948
<< psubstratetap >>
rect 2 15 23 36
rect 33 15 54 36
rect 66 15 87 36
rect 99 15 120 36
rect 132 15 153 36
rect 165 15 186 36
rect 198 15 219 36
rect 231 15 252 36
rect 264 15 285 36
<< nsubstratetap >>
rect 2 1146 23 1167
rect 33 1146 54 1167
rect 66 1146 87 1167
rect 99 1146 120 1167
rect 132 1146 153 1167
rect 165 1146 186 1167
rect 198 1146 219 1167
rect 231 1146 252 1167
rect 264 1146 285 1167
<< metal1 >>
rect 0 1167 291 1176
rect 0 1146 2 1167
rect 23 1146 33 1167
rect 54 1146 66 1167
rect 87 1146 99 1167
rect 120 1146 132 1167
rect 153 1146 165 1167
rect 186 1146 198 1167
rect 219 1146 231 1167
rect 252 1146 264 1167
rect 285 1146 291 1167
rect 11 974 30 1146
rect 114 1110 135 1146
rect 42 974 63 1021
rect 149 1122 265 1134
rect 149 1110 170 1122
rect 78 998 99 1021
rect 78 986 161 998
rect 194 974 215 1021
rect 11 960 215 974
rect 42 948 63 960
rect 194 948 215 960
rect 114 847 135 859
rect 50 826 60 845
rect 114 835 211 847
rect 0 546 291 558
rect 0 517 291 529
rect 0 488 291 500
rect 0 459 291 471
rect 0 430 291 442
rect 78 267 214 279
rect 78 255 99 267
rect 42 194 63 206
rect 114 194 135 206
rect 42 182 135 194
rect 42 158 161 170
rect 42 122 63 158
rect 194 146 215 206
rect 114 134 215 146
rect 114 122 135 134
rect 194 122 215 134
rect 114 36 135 73
rect 149 61 170 73
rect 149 48 265 61
rect 0 15 2 36
rect 23 15 33 36
rect 54 15 66 36
rect 87 15 99 36
rect 120 15 132 36
rect 153 15 165 36
rect 186 15 198 36
rect 219 15 231 36
rect 252 15 264 36
rect 285 15 291 36
rect 0 6 291 15
<< m2contact >>
rect 265 1115 284 1134
rect 231 1086 232 1105
rect 232 1086 250 1105
rect 31 826 50 845
rect 96 800 119 823
rect 231 103 232 122
rect 232 103 250 122
rect 265 48 284 67
<< metal2 >>
rect 33 845 47 1182
rect 33 0 47 826
rect 99 823 113 1182
rect 231 1105 245 1182
rect 264 1134 278 1182
rect 264 1115 265 1134
rect 99 0 113 800
rect 231 122 245 1086
rect 231 0 245 103
rect 264 67 278 1115
rect 264 48 265 67
rect 264 0 278 48
<< labels >>
rlabel metal1 0 6 0 36 3 GND!
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel polysilicon 70 62 70 62 1 A
rlabel metal2 106 62 106 62 1 B
rlabel polysilicon 177 62 177 62 1 nC
rlabel polysilicon 225 62 225 62 1 nS
rlabel metal2 99 0 113 0 1 B
rlabel polysilicon 70 1126 70 1126 1 A
rlabel metal2 106 1126 106 1126 1 B
rlabel polysilicon 224 1121 224 1121 1 nS
rlabel polysilicon 177 1121 177 1121 1 nC
rlabel metal2 99 1182 113 1182 5 B
rlabel metal2 33 1182 47 1182 5 A
rlabel metal2 33 0 47 0 1 A
rlabel metal2 231 1182 245 1182 5 S
rlabel metal2 231 0 245 0 1 S
rlabel metal2 264 0 278 0 1 C
rlabel metal2 264 1182 278 1182 5 C
rlabel metal1 291 1146 291 1176 7 Vdd!
rlabel metal1 291 6 291 36 7 GND!
rlabel metal1 291 546 291 558 7 Scan
rlabel metal1 291 488 291 500 7 Test
rlabel metal1 291 459 291 471 7 Clock
rlabel metal1 291 430 291 442 7 nReset
rlabel metal1 291 517 291 529 7 ScanReturn
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 0 546 0 558 3 Scan
rlabel metal1 0 430 0 442 3 nReset
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 488 0 500 3 Test
<< end >>
