magic
tech tsmc180
timestamp 1733141543
<< nwell >>
rect 0 637 593 1176
<< polysilicon >>
rect 31 1119 40 1131
rect 69 1119 78 1131
rect 31 994 40 1030
rect 69 994 78 1030
rect 105 994 114 1131
rect 141 994 150 1131
rect 31 504 40 905
rect 31 198 40 483
rect 69 198 78 905
rect 105 869 114 905
rect 105 198 114 848
rect 141 563 150 905
rect 179 893 188 1131
rect 179 592 188 872
rect 249 915 258 1141
rect 287 1053 296 1141
rect 325 1110 334 1141
rect 325 1089 329 1110
rect 325 1053 334 1089
rect 363 1053 372 1141
rect 399 1053 408 1141
rect 249 757 258 826
rect 287 757 296 964
rect 325 915 334 964
rect 363 915 372 964
rect 399 915 408 964
rect 141 198 150 542
rect 179 255 188 571
rect 249 352 258 668
rect 287 475 296 668
rect 287 352 296 454
rect 31 112 40 149
rect 69 112 78 149
rect 31 44 40 63
rect 69 44 78 63
rect 105 44 114 149
rect 141 44 150 149
rect 179 44 188 234
rect 249 245 258 303
rect 249 41 258 196
rect 287 147 296 303
rect 325 245 334 826
rect 363 790 372 826
rect 368 769 372 790
rect 363 757 372 769
rect 399 757 408 826
rect 437 814 446 1141
rect 475 1053 484 1141
rect 515 1134 524 1141
rect 515 1053 524 1113
rect 437 757 446 793
rect 363 352 372 668
rect 399 446 408 668
rect 437 562 446 668
rect 475 593 484 964
rect 515 915 524 964
rect 553 915 562 1141
rect 399 352 408 425
rect 437 352 446 541
rect 363 278 372 303
rect 363 245 372 257
rect 399 245 408 303
rect 437 278 446 303
rect 325 147 334 196
rect 363 147 372 196
rect 399 147 408 196
rect 287 41 296 98
rect 325 93 334 98
rect 325 41 334 72
rect 363 41 372 98
rect 399 41 408 98
rect 437 41 446 257
rect 475 147 484 572
rect 515 245 524 826
rect 553 757 562 826
rect 553 591 562 668
rect 553 352 562 570
rect 553 245 562 303
rect 515 147 524 196
rect 475 41 484 98
rect 515 69 524 98
rect 515 41 524 48
rect 553 41 562 196
<< ndiffusion >>
rect 246 303 249 352
rect 258 303 287 352
rect 296 303 299 352
rect 28 149 31 198
rect 40 149 44 198
rect 65 149 69 198
rect 78 149 105 198
rect 114 149 117 198
rect 138 149 141 198
rect 150 149 153 198
rect 28 63 31 112
rect 40 63 43 112
rect 360 303 363 352
rect 372 303 399 352
rect 408 303 437 352
rect 446 303 449 352
rect 322 196 325 245
rect 334 196 363 245
rect 372 196 399 245
rect 408 196 411 245
rect 284 98 287 147
rect 296 98 325 147
rect 334 98 363 147
rect 372 98 399 147
rect 408 98 411 147
rect 512 196 515 245
rect 524 196 553 245
rect 562 196 565 245
rect 472 98 475 147
rect 484 98 515 147
rect 524 98 527 147
<< pdiffusion >>
rect 28 1030 31 1119
rect 40 1030 43 1119
rect 28 905 31 994
rect 40 905 43 994
rect 64 905 69 994
rect 78 905 81 994
rect 102 905 105 994
rect 114 905 117 994
rect 138 905 141 994
rect 150 905 153 994
rect 284 964 287 1053
rect 296 964 299 1053
rect 320 964 325 1053
rect 334 964 337 1053
rect 358 964 363 1053
rect 372 964 375 1053
rect 396 964 399 1053
rect 408 964 411 1053
rect 322 826 325 915
rect 334 826 337 915
rect 358 826 363 915
rect 372 826 375 915
rect 396 826 399 915
rect 408 826 411 915
rect 246 668 249 757
rect 258 668 261 757
rect 282 668 287 757
rect 296 668 299 757
rect 472 964 475 1053
rect 484 964 487 1053
rect 508 964 515 1053
rect 524 964 527 1053
rect 360 668 363 757
rect 372 668 375 757
rect 396 668 399 757
rect 408 668 411 757
rect 432 668 437 757
rect 446 668 449 757
rect 510 826 515 915
rect 524 826 527 915
rect 548 826 553 915
rect 562 826 565 915
<< pohmic >>
rect 0 15 15 36
rect 36 15 101 36
rect 122 15 159 36
rect 180 15 211 36
rect 232 15 263 36
rect 284 15 339 36
rect 360 15 413 36
rect 434 15 487 36
rect 508 15 564 36
rect 585 15 593 36
<< nohmic >>
rect 0 1146 20 1167
rect 41 1146 97 1167
rect 118 1146 162 1167
rect 183 1146 218 1167
rect 239 1146 261 1167
rect 282 1146 339 1167
rect 360 1146 412 1167
rect 433 1146 491 1167
rect 512 1146 563 1167
rect 584 1146 593 1167
<< ntransistor >>
rect 249 303 258 352
rect 287 303 296 352
rect 31 149 40 198
rect 69 149 78 198
rect 105 149 114 198
rect 141 149 150 198
rect 31 63 40 112
rect 363 303 372 352
rect 399 303 408 352
rect 437 303 446 352
rect 325 196 334 245
rect 363 196 372 245
rect 399 196 408 245
rect 287 98 296 147
rect 325 98 334 147
rect 363 98 372 147
rect 399 98 408 147
rect 515 196 524 245
rect 553 196 562 245
rect 475 98 484 147
rect 515 98 524 147
<< ptransistor >>
rect 31 1030 40 1119
rect 31 905 40 994
rect 69 905 78 994
rect 105 905 114 994
rect 141 905 150 994
rect 287 964 296 1053
rect 325 964 334 1053
rect 363 964 372 1053
rect 399 964 408 1053
rect 325 826 334 915
rect 363 826 372 915
rect 399 826 408 915
rect 249 668 258 757
rect 287 668 296 757
rect 475 964 484 1053
rect 515 964 524 1053
rect 363 668 372 757
rect 399 668 408 757
rect 437 668 446 757
rect 515 826 524 915
rect 553 826 562 915
<< polycontact >>
rect 69 1030 90 1119
rect 25 483 46 504
rect 93 848 120 869
rect 167 872 188 893
rect 329 1089 350 1110
rect 249 826 270 915
rect 167 571 188 592
rect 133 542 154 563
rect 287 454 308 475
rect 167 234 188 255
rect 69 63 90 112
rect 249 196 270 245
rect 347 769 368 790
rect 503 1113 524 1134
rect 429 793 450 814
rect 463 572 484 593
rect 425 541 446 562
rect 399 425 420 446
rect 351 257 372 278
rect 431 257 452 278
rect 325 72 346 93
rect 541 668 562 757
rect 548 570 569 591
rect 541 303 562 352
rect 503 48 524 69
<< ndiffcontact >>
rect 225 303 246 352
rect 299 303 320 352
rect 7 149 28 198
rect 44 149 65 198
rect 117 149 138 198
rect 153 149 174 198
rect 7 63 28 112
rect 43 63 64 112
rect 339 303 360 352
rect 449 303 470 352
rect 301 196 322 245
rect 411 196 432 245
rect 263 98 284 147
rect 411 98 432 147
rect 489 196 512 245
rect 565 196 586 245
rect 451 98 472 147
rect 527 98 548 147
<< pdiffcontact >>
rect 7 1030 28 1119
rect 43 1030 64 1119
rect 7 905 28 994
rect 43 905 64 994
rect 81 905 102 994
rect 117 905 138 994
rect 153 905 174 994
rect 263 964 284 1053
rect 299 964 320 1053
rect 337 964 358 1053
rect 375 964 396 1053
rect 411 964 432 1053
rect 301 826 322 915
rect 337 826 358 915
rect 375 826 396 915
rect 411 826 432 915
rect 225 668 246 757
rect 261 668 282 757
rect 299 668 320 757
rect 451 964 472 1053
rect 487 964 508 1053
rect 527 964 548 1053
rect 339 668 360 757
rect 375 668 396 757
rect 411 668 432 757
rect 449 668 470 757
rect 489 826 510 915
rect 527 826 548 915
rect 565 826 586 915
<< psubstratetap >>
rect 15 15 36 36
rect 101 15 122 36
rect 159 15 180 36
rect 211 15 232 36
rect 263 15 284 36
rect 339 15 360 36
rect 413 15 434 36
rect 487 15 508 36
rect 564 15 585 36
<< nsubstratetap >>
rect 20 1146 41 1167
rect 97 1146 118 1167
rect 162 1146 183 1167
rect 218 1146 239 1167
rect 261 1146 282 1167
rect 339 1146 360 1167
rect 412 1146 433 1167
rect 491 1146 512 1167
rect 563 1146 584 1167
<< metal1 >>
rect 0 1167 593 1176
rect 0 1146 20 1167
rect 41 1146 97 1167
rect 118 1146 162 1167
rect 183 1146 218 1167
rect 239 1146 261 1167
rect 282 1146 339 1167
rect 360 1146 412 1167
rect 433 1146 491 1167
rect 512 1146 563 1167
rect 584 1146 593 1167
rect 7 1119 28 1146
rect 64 1030 69 1119
rect 7 994 28 1030
rect 43 1006 138 1018
rect 43 994 64 1006
rect 117 994 138 1006
rect 153 994 174 1146
rect 201 952 231 1146
rect 299 1122 503 1134
rect 299 1077 317 1122
rect 350 1089 508 1101
rect 299 1065 396 1077
rect 299 1053 320 1065
rect 375 1053 396 1065
rect 487 1053 508 1089
rect 263 952 284 964
rect 337 952 358 964
rect 411 952 432 964
rect 451 952 472 964
rect 527 952 548 964
rect 201 927 548 952
rect 86 893 98 905
rect 86 881 167 893
rect 201 757 231 927
rect 337 915 358 927
rect 411 915 432 927
rect 527 915 548 927
rect 270 826 301 915
rect 301 814 322 826
rect 375 814 396 826
rect 489 814 510 826
rect 565 814 586 826
rect 301 802 396 814
rect 450 793 586 814
rect 261 769 347 790
rect 380 769 470 781
rect 261 757 282 769
rect 380 757 396 769
rect 449 757 470 769
rect 201 668 225 757
rect 201 656 246 668
rect 299 656 320 668
rect 470 668 541 757
rect 339 656 360 668
rect 411 656 432 668
rect 201 644 432 656
rect 188 575 463 587
rect 544 571 548 590
rect 0 546 133 558
rect 195 546 425 558
rect 446 546 492 558
rect 511 546 593 558
rect 0 517 593 529
rect 0 488 25 500
rect 46 488 593 500
rect 0 459 287 471
rect 308 459 593 471
rect 0 430 399 442
rect 420 430 593 442
rect 201 364 360 376
rect 201 352 246 364
rect 339 352 360 364
rect 201 303 225 352
rect 470 303 541 352
rect 48 234 167 246
rect 48 198 60 234
rect 87 210 174 222
rect 7 137 28 149
rect 87 137 99 210
rect 153 198 174 210
rect 7 125 99 137
rect 201 184 231 303
rect 299 278 320 303
rect 299 257 351 278
rect 452 257 512 278
rect 489 245 512 257
rect 270 196 301 245
rect 411 184 432 196
rect 565 184 586 196
rect 201 159 586 184
rect 64 63 69 112
rect 7 36 28 63
rect 117 36 138 149
rect 201 36 231 159
rect 411 147 432 159
rect 527 147 548 159
rect 263 60 284 98
rect 451 86 472 98
rect 346 74 472 86
rect 263 48 503 60
rect 0 15 15 36
rect 36 15 101 36
rect 122 15 159 36
rect 180 15 211 36
rect 232 15 263 36
rect 284 15 339 36
rect 360 15 413 36
rect 434 15 487 36
rect 508 15 564 36
rect 585 15 593 36
rect 0 6 593 15
<< m2contact >>
rect 93 848 120 869
rect 525 571 544 590
rect 492 541 511 560
<< metal2 >>
rect 99 869 113 1182
rect 99 0 113 848
rect 495 560 509 1182
rect 528 590 542 1182
rect 495 0 509 541
rect 528 0 542 571
<< labels >>
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel metal1 0 6 0 36 3 GND!
rlabel metal2 99 0 113 0 1 D
rlabel metal2 99 1182 113 1182 5 D
rlabel metal1 593 6 593 36 7 GND!
rlabel metal1 593 517 593 529 7 ScanReturn
rlabel metal1 593 546 593 558 7 Q
rlabel metal1 593 488 593 500 7 Test
rlabel metal1 593 459 593 471 7 Clock
rlabel metal1 593 430 593 442 7 nReset
rlabel metal1 0 430 0 442 3 nReset
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 0 546 0 558 3 SDI
rlabel metal2 495 1182 509 1182 5 Q
rlabel metal2 495 0 509 0 1 Q
rlabel metal2 528 0 542 0 1 nQ
rlabel metal2 528 1182 542 1182 5 nQ
rlabel metal1 593 1146 593 1176 7 Vdd!
<< end >>
