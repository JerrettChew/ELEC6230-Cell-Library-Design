magic
tech tsmc180
timestamp 1733142295
<< nwell >>
rect 0 637 113 1176
<< polysilicon >>
rect 31 1119 40 1130
rect 67 1119 76 1130
rect 31 985 40 1030
rect 67 1018 76 1030
rect 31 112 40 964
rect 67 145 76 997
rect 67 112 76 124
rect 31 52 40 63
rect 67 52 76 63
<< ndiffusion >>
rect 28 63 31 112
rect 40 63 43 112
rect 64 63 67 112
rect 76 63 79 112
<< pdiffusion >>
rect 28 1030 31 1119
rect 40 1030 43 1119
rect 64 1030 67 1119
rect 76 1030 79 1119
<< pohmic >>
rect 0 15 21 36
rect 42 15 63 36
rect 84 15 113 36
<< nohmic >>
rect 0 1146 21 1167
rect 42 1146 63 1167
rect 84 1146 113 1167
<< ntransistor >>
rect 31 63 40 112
rect 67 63 76 112
<< ptransistor >>
rect 31 1030 40 1119
rect 67 1030 76 1119
<< polycontact >>
rect 61 997 82 1018
rect 23 964 44 985
rect 61 124 82 145
<< ndiffcontact >>
rect 7 63 28 112
rect 43 63 64 112
rect 79 63 106 112
<< pdiffcontact >>
rect 7 1030 28 1119
rect 43 1030 64 1119
rect 79 1030 106 1119
<< psubstratetap >>
rect 21 15 42 36
rect 63 15 84 36
<< nsubstratetap >>
rect 21 1146 42 1167
rect 63 1146 84 1167
<< metal1 >>
rect 0 1167 113 1176
rect 0 1146 21 1167
rect 42 1146 63 1167
rect 84 1146 113 1167
rect 43 1119 64 1146
rect 7 1014 19 1030
rect 7 1002 61 1014
rect 94 985 106 1030
rect 82 973 106 985
rect 0 546 113 558
rect 0 517 113 529
rect 0 488 113 500
rect 0 459 113 471
rect 0 430 113 442
rect 83 157 106 169
rect 7 129 61 141
rect 7 112 19 129
rect 94 112 106 157
rect 43 36 64 63
rect 0 15 21 36
rect 42 15 63 36
rect 84 15 113 36
rect 0 6 113 15
<< m2contact >>
rect 30 966 44 985
rect 44 966 49 985
rect 63 966 82 985
rect 64 157 83 176
<< metal2 >>
rect 33 985 47 1182
rect 66 985 80 1182
rect 33 0 47 966
rect 66 176 80 966
rect 66 0 80 157
<< labels >>
rlabel metal1 0 6 0 36 3 GND!
rlabel metal2 66 0 80 0 1 Y
rlabel metal1 113 6 113 36 7 GND!
rlabel metal2 33 0 47 0 1 A
rlabel metal1 0 430 0 442 3 nReset
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 0 546 0 558 3 Scan
rlabel metal1 113 430 113 442 7 nReset
rlabel metal1 113 459 113 471 7 Clock
rlabel metal1 113 488 113 500 7 Test
rlabel metal1 113 517 113 529 7 ScanReturn
rlabel metal1 113 546 113 558 7 Scan
rlabel metal2 66 1182 80 1182 5 Y
rlabel metal2 33 1182 47 1182 5 A
rlabel metal1 113 1146 113 1176 7 Vdd!
rlabel metal1 0 1146 0 1176 3 Vdd!
<< end >>
