magic
tech tsmc180
timestamp 1733141677
<< nwell >>
rect 0 637 391 1176
<< polysilicon >>
rect 31 994 40 1133
rect 142 1119 151 1133
rect 71 994 80 1030
rect 142 994 151 1030
rect 180 994 189 1133
rect 218 1119 227 1133
rect 218 994 227 1030
rect 289 994 298 1133
rect 325 994 334 1030
rect 373 994 382 1134
rect 31 591 40 905
rect 31 200 40 570
rect 71 200 80 905
rect 142 845 151 905
rect 180 845 189 905
rect 142 200 151 824
rect 180 200 189 824
rect 218 504 227 905
rect 289 563 298 905
rect 218 200 227 483
rect 289 200 298 542
rect 325 233 334 905
rect 373 869 382 905
rect 373 592 382 848
rect 373 299 382 571
rect 325 200 334 212
rect 31 44 40 151
rect 71 112 80 151
rect 142 112 151 151
rect 142 44 151 63
rect 180 44 189 151
rect 218 112 227 151
rect 218 44 227 63
rect 289 44 298 151
rect 325 44 334 151
rect 372 44 381 278
<< ndiffusion >>
rect 28 151 31 200
rect 40 151 71 200
rect 80 151 93 200
rect 114 151 142 200
rect 151 151 180 200
rect 189 151 192 200
rect 213 151 218 200
rect 227 151 289 200
rect 298 151 301 200
rect 322 151 325 200
rect 334 151 346 200
rect 139 63 142 112
rect 151 63 154 112
rect 215 63 218 112
rect 227 63 263 112
<< pdiffusion >>
rect 139 1030 142 1119
rect 151 1030 154 1119
rect 215 1030 218 1119
rect 227 1030 263 1119
rect 28 905 31 994
rect 40 905 45 994
rect 66 905 71 994
rect 80 905 83 994
rect 139 905 142 994
rect 151 905 155 994
rect 176 905 180 994
rect 189 905 194 994
rect 215 905 218 994
rect 227 905 230 994
rect 251 905 289 994
rect 298 905 301 994
rect 322 905 325 994
rect 334 905 337 994
<< pohmic >>
rect 0 15 44 36
rect 65 15 99 36
rect 120 15 194 36
rect 215 15 253 36
rect 274 15 301 36
rect 322 15 344 36
rect 365 15 391 36
<< nohmic >>
rect 0 1146 49 1167
rect 70 1146 109 1167
rect 130 1146 185 1167
rect 206 1146 231 1167
rect 252 1146 304 1167
rect 325 1146 360 1167
rect 381 1146 391 1167
<< ntransistor >>
rect 31 151 40 200
rect 71 151 80 200
rect 142 151 151 200
rect 180 151 189 200
rect 218 151 227 200
rect 289 151 298 200
rect 325 151 334 200
rect 142 63 151 112
rect 218 63 227 112
<< ptransistor >>
rect 142 1030 151 1119
rect 218 1030 227 1119
rect 31 905 40 994
rect 71 905 80 994
rect 142 905 151 994
rect 180 905 189 994
rect 218 905 227 994
rect 289 905 298 994
rect 325 905 334 994
<< polycontact >>
rect 71 1030 92 1119
rect 313 1030 334 1119
rect 363 905 384 994
rect 25 570 46 591
rect 132 824 153 845
rect 174 824 195 845
rect 277 542 298 563
rect 212 483 233 504
rect 361 848 382 869
rect 361 571 382 592
rect 361 278 382 299
rect 313 212 334 233
rect 71 63 92 112
<< ndiffcontact >>
rect 7 151 28 200
rect 93 151 114 200
rect 192 151 213 200
rect 301 151 322 200
rect 346 151 367 200
rect 118 63 139 112
rect 154 63 175 112
rect 194 63 215 112
rect 263 63 284 112
<< pdiffcontact >>
rect 118 1030 139 1119
rect 154 1030 175 1119
rect 194 1030 215 1119
rect 263 1030 284 1119
rect 7 905 28 994
rect 45 905 66 994
rect 83 905 104 994
rect 118 905 139 994
rect 155 905 176 994
rect 194 905 215 994
rect 230 905 251 994
rect 301 905 322 994
rect 337 905 358 994
<< psubstratetap >>
rect 44 15 65 36
rect 99 15 120 36
rect 194 15 215 36
rect 253 15 274 36
rect 301 15 322 36
rect 344 15 365 36
<< nsubstratetap >>
rect 49 1146 70 1167
rect 109 1146 130 1167
rect 185 1146 206 1167
rect 231 1146 252 1167
rect 304 1146 325 1167
rect 360 1146 381 1167
<< metal1 >>
rect 0 1167 391 1176
rect 0 1146 49 1167
rect 70 1146 109 1167
rect 130 1146 185 1167
rect 206 1146 231 1167
rect 252 1146 304 1167
rect 325 1146 360 1167
rect 381 1146 391 1167
rect 154 1119 175 1146
rect 92 1030 118 1119
rect 194 1119 215 1146
rect 7 1006 104 1018
rect 7 994 28 1006
rect 83 994 104 1006
rect 45 869 66 905
rect 118 1006 215 1018
rect 118 994 139 1006
rect 194 994 215 1006
rect 230 994 251 1146
rect 284 1030 313 1119
rect 358 905 363 994
rect 83 893 104 905
rect 155 893 175 905
rect 83 881 175 893
rect 194 893 215 905
rect 301 893 322 905
rect 194 881 322 893
rect 45 857 361 869
rect 46 575 322 587
rect 0 546 277 558
rect 310 558 322 575
rect 382 575 391 587
rect 310 546 391 558
rect 0 517 391 529
rect 0 488 212 500
rect 233 488 391 500
rect 0 459 391 471
rect 0 430 391 442
rect 7 278 361 290
rect 7 200 28 278
rect 93 245 367 266
rect 93 200 114 245
rect 263 214 313 231
rect 7 139 28 151
rect 192 139 213 151
rect 7 124 213 139
rect 263 112 284 214
rect 346 200 367 245
rect 92 63 118 112
rect 154 36 175 63
rect 194 36 215 63
rect 301 36 322 151
rect 0 15 44 36
rect 65 15 99 36
rect 120 15 194 36
rect 215 15 253 36
rect 274 15 301 36
rect 322 15 344 36
rect 365 15 391 36
rect 0 6 391 15
<< m2contact >>
rect 124 824 132 845
rect 132 824 143 845
rect 165 824 174 845
rect 174 824 184 845
<< metal2 >>
rect 132 845 146 1182
rect 143 824 146 845
rect 132 0 146 824
rect 165 845 179 1182
rect 165 0 179 824
<< labels >>
rlabel metal2 132 1182 146 1182 5 Load
rlabel metal2 165 1182 179 1182 5 D
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel metal1 391 1146 391 1176 7 Vdd!
rlabel metal1 391 459 391 471 7 Clock
rlabel metal1 391 488 391 500 7 Test
rlabel metal1 391 517 391 529 7 ScanReturn
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 0 546 0 558 3 SDI
rlabel metal1 391 546 391 558 7 Q
rlabel metal1 0 430 0 442 3 nReset
rlabel metal1 391 430 391 442 7 nReset
rlabel metal1 391 575 391 587 7 nD
rlabel metal2 165 0 179 0 1 D
rlabel metal2 132 0 146 0 1 Load
rlabel metal1 391 6 391 36 7 GND!
rlabel metal1 0 6 0 36 3 GND!
<< end >>
