magic
tech tsmc180
timestamp 1733141893
<< nwell >>
rect 0 637 87 1176
<< polysilicon >>
rect 31 1119 40 1130
rect 31 1018 40 1030
rect 31 112 40 997
rect 31 52 40 63
<< ndiffusion >>
rect 28 63 31 112
rect 40 63 43 112
<< pdiffusion >>
rect 28 1030 31 1119
rect 40 1030 43 1119
<< pohmic >>
rect 0 15 46 36
rect 67 15 87 36
<< nohmic >>
rect 0 1146 46 1167
rect 67 1146 87 1167
<< ntransistor >>
rect 31 63 40 112
<< ptransistor >>
rect 31 1030 40 1119
<< polycontact >>
rect 24 997 45 1018
<< ndiffcontact >>
rect 7 63 28 112
rect 43 63 64 112
<< pdiffcontact >>
rect 7 1030 28 1119
rect 43 1030 64 1119
<< psubstratetap >>
rect 46 15 67 36
<< nsubstratetap >>
rect 46 1146 67 1167
<< metal1 >>
rect 0 1167 87 1176
rect 0 1146 46 1167
rect 67 1146 87 1167
rect 7 1119 28 1146
rect 0 546 87 558
rect 0 517 87 529
rect 0 488 87 500
rect 0 459 87 471
rect 0 430 87 442
rect 7 36 28 63
rect 0 15 46 36
rect 67 15 87 36
rect 0 6 87 15
<< m2contact >>
rect 61 1100 64 1119
rect 64 1100 80 1119
rect 31 999 45 1018
rect 45 999 50 1018
rect 61 63 64 82
rect 64 63 80 82
<< metal2 >>
rect 33 1018 47 1182
rect 66 1119 80 1182
rect 33 0 47 999
rect 66 82 80 1100
rect 66 0 80 63
<< labels >>
rlabel metal2 33 0 47 0 1 A
rlabel metal2 66 0 80 0 1 Y
rlabel metal1 0 6 0 36 3 GND!
rlabel metal1 87 6 87 36 7 GND!
rlabel metal1 0 546 0 558 3 Scan
rlabel metal1 0 517 0 529 3 ScanReturn
rlabel metal1 0 488 0 500 3 Test
rlabel metal1 0 459 0 471 3 Clock
rlabel metal1 0 430 0 442 3 nReset
rlabel metal1 87 546 87 558 7 Scan
rlabel metal1 87 517 87 529 7 ScanReturn
rlabel metal1 87 488 87 500 7 Test
rlabel metal1 87 459 87 471 7 Clock
rlabel metal1 87 430 87 442 7 nReset
rlabel metal1 87 1146 87 1176 7 Vdd!
rlabel metal1 0 1146 0 1176 3 Vdd!
rlabel metal2 66 1182 80 1182 5 Y
rlabel metal2 33 1182 47 1182 5 A
<< end >>
